`timescale 1 ns/100 ps
// Version: v11.8 11.8.0.26


module MSS_005(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module u8_sb_HPMS(
       CoreAHBLite_0_AHBmslave16_HWDATA,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0,
       CoreAHBLite_0_AHBmslave16_HTRANS_0,
       CoreAHBLite_0_AHBmslave16_HSIZE_0,
       CoreAHBLite_0_AHBmslave16_HADDR_0,
       CoreAHBLite_0_AHBmslave16_HADDR_1,
       CoreAHBLite_0_AHBmslave16_HADDR_2,
       CoreAHBLite_0_AHBmslave16_HADDR_3,
       CoreAHBLite_0_AHBmslave16_HADDR_4,
       CoreAHBLite_0_AHBmslave16_HADDR_5,
       CoreAHBLite_0_AHBmslave16_HADDR_6,
       CoreAHBLite_0_AHBmslave16_HADDR_7,
       CoreAHBLite_0_AHBmslave16_HADDR_8,
       CoreAHBLite_0_AHBmslave16_HADDR_9,
       CoreAHBLite_0_AHBmslave16_HADDR_10,
       CoreAHBLite_0_AHBmslave16_HADDR_11,
       CoreAHBLite_0_AHBmslave16_HADDR_12,
       CoreAHBLite_0_AHBmslave16_HADDR_13,
       CoreAHBLite_0_AHBmslave16_HADDR_14,
       CoreAHBLite_0_AHBmslave16_HADDR_27,
       CoreAHBLite_0_AHBmslave16_HADDR_28,
       masterAddrInProg_0,
       GL0_INST,
       u8_sb_0_FIC_0_LOCK,
       CoreAHBLite_0_AHBmslave16_HWRITE,
       N_128_i,
       u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F,
       u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N,
       m0s16DataSel,
       CoreAHBLite_0_AHBmslave16_HREADY_m_0,
       CoreAHBLite_0_AHBmslave16_HREADY
    );
input  [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
output [31:0] u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0;
input  CoreAHBLite_0_AHBmslave16_HTRANS_0;
input  CoreAHBLite_0_AHBmslave16_HSIZE_0;
input  CoreAHBLite_0_AHBmslave16_HADDR_0;
input  CoreAHBLite_0_AHBmslave16_HADDR_1;
input  CoreAHBLite_0_AHBmslave16_HADDR_2;
input  CoreAHBLite_0_AHBmslave16_HADDR_3;
input  CoreAHBLite_0_AHBmslave16_HADDR_4;
input  CoreAHBLite_0_AHBmslave16_HADDR_5;
input  CoreAHBLite_0_AHBmslave16_HADDR_6;
input  CoreAHBLite_0_AHBmslave16_HADDR_7;
input  CoreAHBLite_0_AHBmslave16_HADDR_8;
input  CoreAHBLite_0_AHBmslave16_HADDR_9;
input  CoreAHBLite_0_AHBmslave16_HADDR_10;
input  CoreAHBLite_0_AHBmslave16_HADDR_11;
input  CoreAHBLite_0_AHBmslave16_HADDR_12;
input  CoreAHBLite_0_AHBmslave16_HADDR_13;
input  CoreAHBLite_0_AHBmslave16_HADDR_14;
input  CoreAHBLite_0_AHBmslave16_HADDR_27;
input  CoreAHBLite_0_AHBmslave16_HADDR_28;
input  masterAddrInProg_0;
input  GL0_INST;
input  u8_sb_0_FIC_0_LOCK;
input  CoreAHBLite_0_AHBmslave16_HWRITE;
input  N_128_i;
output u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F;
output u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N;
input  m0s16DataSel;
output CoreAHBLite_0_AHBmslave16_HREADY_m_0;
inout  CoreAHBLite_0_AHBmslave16_HREADY;

    wire \CoreAHBLite_0_AHBmslave16_HRDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[0] , VCC_net_1, GND_net_1;
    
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_6 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[7] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_0 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[1] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_24 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[25] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_14 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[15] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_23 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[24] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_13 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[14] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14]));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_4 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[5] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_29 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[30] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_19 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[20] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_7 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[8] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8]));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_30 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[31] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_3 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[4] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_26 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[27] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_20 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[21] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21]));
    MSS_005 #( .INIT(1438'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C00000000609300000003FFFFE000000000000010000000000F15C000001FE5FE4010842108421000001FE34001FF8000000000000000020051127FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(49.152)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({\CoreAHBLite_0_AHBmslave16_HRDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[0] }), .F_FM0_READYOUT(
        CoreAHBLite_0_AHBmslave16_HREADY), .F_FM0_RESP(), .F_HM0_ADDR({
        nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17, nc18, 
        nc19, nc20, nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, 
        nc29, nc30, nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, 
        nc39}), .F_HM0_ENABLE(), .F_HM0_SEL(), .F_HM0_SIZE({nc40, nc41})
        , .F_HM0_TRANS1(), .F_HM0_WDATA({nc42, nc43, nc44, nc45, nc46, 
        nc47, nc48, nc49, nc50, nc51, nc52, nc53, nc54, nc55, nc56, 
        nc57, nc58, nc59, nc60, nc61, nc62, nc63, nc64, nc65, nc66, 
        nc67, nc68, nc69, nc70, nc71, nc72, nc73}), .F_HM0_WRITE(), 
        .FAB_CHRGVBUS(), .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), 
        .FAB_DPPULLDOWN(), .FAB_DRVVBUS(), .FAB_IDPULLUP(), 
        .FAB_OPMODE({nc74, nc75}), .FAB_SUSPENDM(), .FAB_TERMSEL(), 
        .FAB_TXVALID(), .FAB_VCONTROL({nc76, nc77, nc78, nc79}), 
        .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({nc80, nc81}), 
        .FAB_XDATAOUT({nc82, nc83, nc84, nc85, nc86, nc87, nc88, nc89})
        , .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc90, nc91}), 
        .FIC32_1_MASTER({nc92, nc93}), .FPGA_RESET_N(
        u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F), .GTX_CLK(), .H2F_INTERRUPT({
        nc94, nc95, nc96, nc97, nc98, nc99, nc100, nc101, nc102, nc103, 
        nc104, nc105, nc106, nc107, nc108, nc109}), .H2F_NMI(), 
        .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc110, nc111, nc112, nc113, nc114, nc115, 
        nc116, nc117, nc118, nc119, nc120, nc121, nc122, nc123}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc124, nc125, nc126, nc127, nc128, nc129, 
        nc130, nc131, nc132, nc133, nc134, nc135, nc136, nc137, nc138, 
        nc139, nc140, nc141, nc142, nc143, nc144, nc145, nc146, nc147, 
        nc148, nc149, nc150, nc151, nc152, nc153, nc154, nc155}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc156, nc157, nc158, nc159, 
        nc160, nc161, nc162, nc163, nc164, nc165}), .TRACECLK(), 
        .TRACEDATA({nc166, nc167, nc168, nc169}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc170, nc171, nc172, 
        nc173}), .TXDF({nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc182, nc183, nc184, nc185})
        , .F_BRESP_HRESP0({nc186, nc187}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc188, nc189, nc190, nc191, nc192, nc193, 
        nc194, nc195, nc196, nc197, nc198, nc199, nc200, nc201, nc202, 
        nc203, nc204, nc205, nc206, nc207, nc208, nc209, nc210, nc211, 
        nc212, nc213, nc214, nc215, nc216, nc217, nc218, nc219, nc220, 
        nc221, nc222, nc223, nc224, nc225, nc226, nc227, nc228, nc229, 
        nc230, nc231, nc232, nc233, nc234, nc235, nc236, nc237, nc238, 
        nc239, nc240, nc241, nc242, nc243, nc244, nc245, nc246, nc247, 
        nc248, nc249, nc250, nc251}), .F_RID({nc252, nc253, nc254, 
        nc255}), .F_RLAST(), .F_RRESP_HRESP1({nc256, nc257}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc258, nc259, 
        nc260, nc261, nc262, nc263, nc264, nc265, nc266, nc267, nc268, 
        nc269, nc270, nc271, nc272, nc273}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F2HCALIB(VCC_net_1), 
        .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({GND_net_1, 
        CoreAHBLite_0_AHBmslave16_HADDR_28, 
        CoreAHBLite_0_AHBmslave16_HADDR_27, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        CoreAHBLite_0_AHBmslave16_HADDR_14, 
        CoreAHBLite_0_AHBmslave16_HADDR_14, 
        CoreAHBLite_0_AHBmslave16_HADDR_13, 
        CoreAHBLite_0_AHBmslave16_HADDR_12, 
        CoreAHBLite_0_AHBmslave16_HADDR_11, 
        CoreAHBLite_0_AHBmslave16_HADDR_10, 
        CoreAHBLite_0_AHBmslave16_HADDR_9, 
        CoreAHBLite_0_AHBmslave16_HADDR_8, 
        CoreAHBLite_0_AHBmslave16_HADDR_7, 
        CoreAHBLite_0_AHBmslave16_HADDR_6, 
        CoreAHBLite_0_AHBmslave16_HADDR_5, 
        CoreAHBLite_0_AHBmslave16_HADDR_4, 
        CoreAHBLite_0_AHBmslave16_HADDR_3, 
        CoreAHBLite_0_AHBmslave16_HADDR_2, 
        CoreAHBLite_0_AHBmslave16_HADDR_1, 
        CoreAHBLite_0_AHBmslave16_HADDR_0, GND_net_1, GND_net_1}), 
        .F_FM0_ENABLE(GND_net_1), .F_FM0_MASTLOCK(
        CoreAHBLite_0_AHBmslave16_HSIZE_0), .F_FM0_READY(
        CoreAHBLite_0_AHBmslave16_HREADY), .F_FM0_SEL(N_128_i), 
        .F_FM0_SIZE({CoreAHBLite_0_AHBmslave16_HSIZE_0, GND_net_1}), 
        .F_FM0_TRANS1(CoreAHBLite_0_AHBmslave16_HTRANS_0), 
        .F_FM0_WDATA({CoreAHBLite_0_AHBmslave16_HWDATA[31], 
        CoreAHBLite_0_AHBmslave16_HWDATA[30], 
        CoreAHBLite_0_AHBmslave16_HWDATA[29], 
        CoreAHBLite_0_AHBmslave16_HWDATA[28], 
        CoreAHBLite_0_AHBmslave16_HWDATA[27], 
        CoreAHBLite_0_AHBmslave16_HWDATA[26], 
        CoreAHBLite_0_AHBmslave16_HWDATA[25], 
        CoreAHBLite_0_AHBmslave16_HWDATA[24], 
        CoreAHBLite_0_AHBmslave16_HWDATA[23], 
        CoreAHBLite_0_AHBmslave16_HWDATA[22], 
        CoreAHBLite_0_AHBmslave16_HWDATA[21], 
        CoreAHBLite_0_AHBmslave16_HWDATA[20], 
        CoreAHBLite_0_AHBmslave16_HWDATA[19], 
        CoreAHBLite_0_AHBmslave16_HWDATA[18], 
        CoreAHBLite_0_AHBmslave16_HWDATA[17], 
        CoreAHBLite_0_AHBmslave16_HWDATA[16], 
        CoreAHBLite_0_AHBmslave16_HWDATA[15], 
        CoreAHBLite_0_AHBmslave16_HWDATA[14], 
        CoreAHBLite_0_AHBmslave16_HWDATA[13], 
        CoreAHBLite_0_AHBmslave16_HWDATA[12], 
        CoreAHBLite_0_AHBmslave16_HWDATA[11], 
        CoreAHBLite_0_AHBmslave16_HWDATA[10], 
        CoreAHBLite_0_AHBmslave16_HWDATA[9], 
        CoreAHBLite_0_AHBmslave16_HWDATA[8], 
        CoreAHBLite_0_AHBmslave16_HWDATA[7], 
        CoreAHBLite_0_AHBmslave16_HWDATA[6], 
        CoreAHBLite_0_AHBmslave16_HWDATA[5], 
        CoreAHBLite_0_AHBmslave16_HWDATA[4], 
        CoreAHBLite_0_AHBmslave16_HWDATA[3], 
        CoreAHBLite_0_AHBmslave16_HWDATA[2], 
        CoreAHBLite_0_AHBmslave16_HWDATA[1], 
        CoreAHBLite_0_AHBmslave16_HWDATA[0]}), .F_FM0_WRITE(
        CoreAHBLite_0_AHBmslave16_HWRITE), .F_HM0_RDATA({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_HM0_READY(VCC_net_1), .F_HM0_RESP(GND_net_1), 
        .FAB_AVALID(VCC_net_1), .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(
        VCC_net_1), .FAB_LINESTATE({VCC_net_1, VCC_net_1}), 
        .FAB_M3_RESET_N(GND_net_1), .FAB_PLL_LOCK(u8_sb_0_FIC_0_LOCK), 
        .FAB_RXACTIVE(VCC_net_1), .FAB_RXERROR(VCC_net_1), 
        .FAB_RXVALID(VCC_net_1), .FAB_RXVALIDH(GND_net_1), 
        .FAB_SESSEND(VCC_net_1), .FAB_TXREADY(VCC_net_1), 
        .FAB_VBUSVALID(VCC_net_1), .FAB_VSTATUS({VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .FAB_XDATAIN({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .GTX_CLKPF(VCC_net_1), .I2C0_BCLK(VCC_net_1), 
        .I2C0_SCL_F2H_SCP(VCC_net_1), .I2C0_SDA_F2H_SCP(VCC_net_1), 
        .I2C1_BCLK(VCC_net_1), .I2C1_SCL_F2H_SCP(VCC_net_1), 
        .I2C1_SDA_F2H_SCP(VCC_net_1), .MDIF(VCC_net_1), 
        .MGPIO0A_F2H_GPIN(VCC_net_1), .MGPIO10A_F2H_GPIN(VCC_net_1), 
        .MGPIO11A_F2H_GPIN(VCC_net_1), .MGPIO11B_F2H_GPIN(VCC_net_1), 
        .MGPIO12A_F2H_GPIN(VCC_net_1), .MGPIO13A_F2H_GPIN(VCC_net_1), 
        .MGPIO14A_F2H_GPIN(VCC_net_1), .MGPIO15A_F2H_GPIN(VCC_net_1), 
        .MGPIO16A_F2H_GPIN(VCC_net_1), .MGPIO17B_F2H_GPIN(VCC_net_1), 
        .MGPIO18B_F2H_GPIN(VCC_net_1), .MGPIO19B_F2H_GPIN(VCC_net_1), 
        .MGPIO1A_F2H_GPIN(VCC_net_1), .MGPIO20B_F2H_GPIN(VCC_net_1), 
        .MGPIO21B_F2H_GPIN(VCC_net_1), .MGPIO22B_F2H_GPIN(VCC_net_1), 
        .MGPIO24B_F2H_GPIN(VCC_net_1), .MGPIO25B_F2H_GPIN(VCC_net_1), 
        .MGPIO26B_F2H_GPIN(VCC_net_1), .MGPIO27B_F2H_GPIN(VCC_net_1), 
        .MGPIO28B_F2H_GPIN(VCC_net_1), .MGPIO29B_F2H_GPIN(VCC_net_1), 
        .MGPIO2A_F2H_GPIN(VCC_net_1), .MGPIO30B_F2H_GPIN(VCC_net_1), 
        .MGPIO31B_F2H_GPIN(VCC_net_1), .MGPIO3A_F2H_GPIN(VCC_net_1), 
        .MGPIO4A_F2H_GPIN(VCC_net_1), .MGPIO5A_F2H_GPIN(VCC_net_1), 
        .MGPIO6A_F2H_GPIN(VCC_net_1), .MGPIO7A_F2H_GPIN(VCC_net_1), 
        .MGPIO8A_F2H_GPIN(VCC_net_1), .MGPIO9A_F2H_GPIN(VCC_net_1), 
        .MMUART0_CTS_F2H_SCP(VCC_net_1), .MMUART0_DCD_F2H_SCP(
        VCC_net_1), .MMUART0_DSR_F2H_SCP(VCC_net_1), 
        .MMUART0_DTR_F2H_SCP(VCC_net_1), .MMUART0_RI_F2H_SCP(VCC_net_1)
        , .MMUART0_RTS_F2H_SCP(VCC_net_1), .MMUART0_RXD_F2H_SCP(
        VCC_net_1), .MMUART0_SCK_F2H_SCP(VCC_net_1), 
        .MMUART0_TXD_F2H_SCP(VCC_net_1), .MMUART1_CTS_F2H_SCP(
        VCC_net_1), .MMUART1_DCD_F2H_SCP(VCC_net_1), 
        .MMUART1_DSR_F2H_SCP(VCC_net_1), .MMUART1_RI_F2H_SCP(VCC_net_1)
        , .MMUART1_RTS_F2H_SCP(VCC_net_1), .MMUART1_RXD_F2H_SCP(
        VCC_net_1), .MMUART1_SCK_F2H_SCP(VCC_net_1), 
        .MMUART1_TXD_F2H_SCP(VCC_net_1), .PER2_FABRIC_PRDATA({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .PER2_FABRIC_PREADY(VCC_net_1), 
        .PER2_FABRIC_PSLVERR(GND_net_1), .RCGF({VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .RX_CLKPF(VCC_net_1), 
        .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), .RX_EV(VCC_net_1), 
        .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .SLEEPHOLDREQ(GND_net_1), 
        .SMBALERT_NI0(VCC_net_1), .SMBALERT_NI1(VCC_net_1), 
        .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(VCC_net_1), .SPI0_CLK_IN(
        VCC_net_1), .SPI0_SDI_F2H_SCP(VCC_net_1), .SPI0_SDO_F2H_SCP(
        VCC_net_1), .SPI0_SS0_F2H_SCP(VCC_net_1), .SPI0_SS1_F2H_SCP(
        VCC_net_1), .SPI0_SS2_F2H_SCP(VCC_net_1), .SPI0_SS3_F2H_SCP(
        VCC_net_1), .SPI1_CLK_IN(VCC_net_1), .SPI1_SDI_F2H_SCP(
        VCC_net_1), .SPI1_SDO_F2H_SCP(VCC_net_1), .SPI1_SS0_F2H_SCP(
        VCC_net_1), .SPI1_SS1_F2H_SCP(VCC_net_1), .SPI1_SS2_F2H_SCP(
        VCC_net_1), .SPI1_SS3_F2H_SCP(VCC_net_1), .TX_CLKPF(VCC_net_1), 
        .USER_MSS_GPIO_RESET_N(VCC_net_1), .USER_MSS_RESET_N(VCC_net_1)
        , .XCLK_FAB(VCC_net_1), .CLK_BASE(GL0_INST), .CLK_MDDR_APB(
        VCC_net_1), .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .F_ARBURST_HTRANS1({GND_net_1, GND_net_1}), .F_ARID_HSEL1({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_ARLOCK_HMASTLOCK1({GND_net_1, GND_net_1}), .F_ARSIZE_HSIZE1({
        GND_net_1, GND_net_1}), .F_ARVALID_HWRITE1(GND_net_1), 
        .F_AWADDR_HADDR0({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_AWBURST_HTRANS0({
        GND_net_1, GND_net_1}), .F_AWID_HSEL0({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_AWLEN_HBURST0({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_AWLOCK_HMASTLOCK0({GND_net_1, 
        GND_net_1}), .F_AWSIZE_HSIZE0({GND_net_1, GND_net_1}), 
        .F_AWVALID_HWRITE0(GND_net_1), .F_BREADY(GND_net_1), 
        .F_RMW_AXI(GND_net_1), .F_RREADY(GND_net_1), .F_WDATA_HWDATA01({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .F_WID_HREADY01({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .F_WLAST(
        GND_net_1), .F_WSTRB({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_WVALID(GND_net_1), .FPGA_MDDR_ARESET_N(VCC_net_1), 
        .MDDR_FABRIC_PADDR({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .MDDR_FABRIC_PENABLE(VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), 
        .MDDR_FABRIC_PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PWRITE(
        VCC_net_1), .PRESET_N(GND_net_1), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND_net_1), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), .USBC_XCLK_IN(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc274, nc275, 
        nc276, nc277, nc278, nc279, nc280, nc281, nc282, nc283, nc284, 
        nc285, nc286, nc287, nc288, nc289}), .DRAM_BA({nc290, nc291, 
        nc292}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc293, nc294, nc295}), .DRAM_DQ_OUT({nc296, 
        nc297, nc298, nc299, nc300, nc301, nc302, nc303, nc304, nc305, 
        nc306, nc307, nc308, nc309, nc310, nc311, nc312, nc313}), 
        .DRAM_DQS_OUT({nc314, nc315, nc316}), .DRAM_FIFO_WE_OUT({nc317, 
        nc318}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), .USBC_XCLK_OUT(), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc319, nc320, 
        nc321}), .DRAM_DQ_OE({nc322, nc323, nc324, nc325, nc326, nc327, 
        nc328, nc329, nc330, nc331, nc332, nc333, nc334, nc335, nc336, 
        nc337, nc338, nc339}), .DRAM_DQS_OE({nc340, nc341, nc342}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), .USBC_XCLK_OE());
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNIBVGL (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_16 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[17] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_10 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[11] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_21 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[22] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_9 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[10] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_22 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[23] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_11 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[12] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_12 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[13] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[0] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_2 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[3] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_1 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[2] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_8 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[9] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_28 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[29] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_5 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[6] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_18 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[19] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_27 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[28] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_25 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[26] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_17 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[18] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18]));
    CFG2 #( .INIT(4'h8) )  MSS_ADLIB_INST_RNI9FUD_15 (.A(m0s16DataSel), 
        .B(\CoreAHBLite_0_AHBmslave16_HRDATA[16] ), .Y(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16]));
    
endmodule


module CoreResetP_Z5(
       u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N,
       u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F,
       SYSRESET_POR,
       GL0_INST,
       u8_sb_0_HPMS_READY
    );
input  u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N;
input  u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F;
input  SYSRESET_POR;
input  GL0_INST;
output u8_sb_0_HPMS_READY;

    wire MSS_HPMS_READY_int_net_1, mss_ready_select_net_1, VCC_net_1, 
        POWER_ON_RESET_N_clk_base_net_1, mss_ready_select4_net_1, 
        GND_net_1, mss_ready_state_net_1, RESET_N_M2F_clk_base_net_1, 
        POWER_ON_RESET_N_q1_net_1, RESET_N_M2F_q1_net_1, 
        FIC_2_APB_M_PRESET_N_clk_base_net_1, 
        FIC_2_APB_M_PRESET_N_q1_net_1, MSS_HPMS_READY_int_4_net_1;
    
    SLE RESET_N_M2F_clk_base (.D(RESET_N_M2F_q1_net_1), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(RESET_N_M2F_clk_base_net_1));
    SLE POWER_ON_RESET_N_clk_base (.D(POWER_ON_RESET_N_q1_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_clk_base_net_1));
    SLE mss_ready_select (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        mss_ready_select4_net_1), .ALn(POWER_ON_RESET_N_clk_base_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(mss_ready_select_net_1));
    GND GND (.Y(GND_net_1));
    SLE mss_ready_state (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        RESET_N_M2F_clk_base_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_state_net_1));
    CLKINT MSS_HPMS_READY_int_RNIVGLD (.A(MSS_HPMS_READY_int_net_1), 
        .Y(u8_sb_0_HPMS_READY));
    VCC VCC (.Y(VCC_net_1));
    SLE RESET_N_M2F_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_q1_net_1));
    SLE FIC_2_APB_M_PRESET_N_clk_base (.D(
        FIC_2_APB_M_PRESET_N_q1_net_1), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FIC_2_APB_M_PRESET_N_clk_base_net_1));
    SLE POWER_ON_RESET_N_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_q1_net_1));
    CFG2 #( .INIT(4'h8) )  mss_ready_select4 (.A(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .B(mss_ready_state_net_1)
        , .Y(mss_ready_select4_net_1));
    CFG3 #( .INIT(8'hE0) )  MSS_HPMS_READY_int_4 (.A(
        RESET_N_M2F_clk_base_net_1), .B(mss_ready_select_net_1), .C(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .Y(
        MSS_HPMS_READY_int_4_net_1));
    SLE FIC_2_APB_M_PRESET_N_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(FIC_2_APB_M_PRESET_N_q1_net_1));
    SLE MSS_HPMS_READY_int (.D(MSS_HPMS_READY_int_4_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        MSS_HPMS_READY_int_net_1));
    
endmodule


module COREAHBLITE_MASTERSTAGE_1_1_85_65536_0s_0_1_0(
       test_0_HADDR,
       regHADDR,
       masterDataInProg_0,
       M0GATEDHADDR_0,
       M0GATEDHADDR_13,
       test_0_HTRANS_0,
       M0GATEDHSIZE_0,
       test_0_HADDR_i_0,
       CoreAHBLite_0_AHBmslave16_HREADY_m_0,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       CoreAHBLite_0_AHBmslave16_HREADY,
       m0s16AddrSel,
       VCC_0,
       VCC_0_reto,
       d_masterRegAddrSel,
       masterRegAddrSel,
       test_0_HWRITE,
       regHWRITE,
       m0s16DataSel,
       GL0_INST,
       u8_sb_0_HPMS_READY
    );
input  [16:2] test_0_HADDR;
output [15:2] regHADDR;
input  masterDataInProg_0;
output M0GATEDHADDR_0;
output M0GATEDHADDR_13;
input  test_0_HTRANS_0;
output M0GATEDHSIZE_0;
input  test_0_HADDR_i_0;
input  CoreAHBLite_0_AHBmslave16_HREADY_m_0;
output u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
input  CoreAHBLite_0_AHBmslave16_HREADY;
output m0s16AddrSel;
output VCC_0;
input  VCC_0_reto;
output d_masterRegAddrSel;
output masterRegAddrSel;
input  test_0_HWRITE;
output regHWRITE;
output m0s16DataSel;
input  GL0_INST;
input  u8_sb_0_HPMS_READY;

    wire \regHADDR[29]_net_1 , VCC_net_1, masterAddrClockEnable_net_1, 
        GND_net_1, SDATASELInt_54_net_1, \regHADDR[16]_net_1 , 
        regHTRANS_net_1, masterAddrClockEnable4_1_net_1;
    
    CFG3 #( .INIT(8'h8F) )  HREADY_M_0_iv (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(masterDataInProg_0), .C(
        m0s16DataSel), .Y(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0));
    SLE \regHADDR[2]  (.D(test_0_HADDR[2]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[2]));
    SLE \regHADDR[29]  (.D(test_0_HADDR_i_0), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\regHADDR[29]_net_1 ));
    SLE \regHADDR[12]  (.D(test_0_HADDR[12]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[12]));
    CFG4 #( .INIT(16'h0400) )  masterAddrClockEnable (.A(
        masterRegAddrSel), .B(m0s16AddrSel), .C(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0), .D(
        masterAddrClockEnable4_1_net_1), .Y(
        masterAddrClockEnable_net_1));
    SLE regHTRANS (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHTRANS_net_1));
    SLE \regHADDR[13]  (.D(test_0_HADDR[13]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[13]));
    SLE \regHADDR[7]  (.D(test_0_HADDR[7]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[7]));
    SLE \regHADDR[14]  (.D(test_0_HADDR[14]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[14]));
    CFG4 #( .INIT(16'h0C08) )  d_masterRegAddrSel_inst_1 (.A(
        masterRegAddrSel), .B(m0s16AddrSel), .C(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0), .D(
        masterAddrClockEnable4_1_net_1), .Y(d_masterRegAddrSel));
    SLE \regHADDR[4]  (.D(test_0_HADDR[4]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[4]));
    CFG3 #( .INIT(8'hE4) )  GATEDHTRANS (.A(masterRegAddrSel), .B(
        test_0_HTRANS_0), .C(regHTRANS_net_1), .Y(m0s16AddrSel));
    CFG4 #( .INIT(16'h8A0A) )  masterAddrClockEnable4_1 (.A(
        test_0_HTRANS_0), .B(masterDataInProg_0), .C(m0s16DataSel), .D(
        CoreAHBLite_0_AHBmslave16_HREADY), .Y(
        masterAddrClockEnable4_1_net_1));
    GND GND (.Y(GND_net_1));
    SLE \regHADDR[5]  (.D(test_0_HADDR[5]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[5]));
    CFG3 #( .INIT(8'hBA) )  SDATASELInt_54 (.A(m0s16AddrSel), .B(
        CoreAHBLite_0_AHBmslave16_HREADY), .C(m0s16DataSel), .Y(
        SDATASELInt_54_net_1));
    SLE \SDATASELInt[16]  (.D(SDATASELInt_54_net_1), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        m0s16DataSel));
    CFG2 #( .INIT(4'hE) )  regHTRANS_reten (.A(
        masterAddrClockEnable_net_1), .B(VCC_0_reto), .Y(VCC_0));
    CFG3 #( .INIT(8'hB1) )  \PREGATEDHADDR[29]  (.A(masterRegAddrSel), 
        .B(test_0_HADDR[16]), .C(\regHADDR[29]_net_1 ), .Y(
        M0GATEDHADDR_13));
    SLE masterRegAddrSel_inst_1 (.D(d_masterRegAddrSel), .CLK(GL0_INST)
        , .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        masterRegAddrSel));
    CFG3 #( .INIT(8'hE4) )  \PREGATEDHADDR[16]  (.A(masterRegAddrSel), 
        .B(test_0_HADDR[16]), .C(\regHADDR[16]_net_1 ), .Y(
        M0GATEDHADDR_0));
    SLE \regHADDR[11]  (.D(test_0_HADDR[11]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[11]));
    CFG2 #( .INIT(4'hD) )  \GATEDHSIZE[1]  (.A(masterRegAddrSel), .B(
        regHTRANS_net_1), .Y(M0GATEDHSIZE_0));
    SLE regHWRITE_inst_1 (.D(test_0_HWRITE), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHWRITE));
    SLE \regHADDR[3]  (.D(test_0_HADDR[3]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[3]));
    SLE \regHADDR[16]  (.D(test_0_HADDR[16]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\regHADDR[16]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \regHADDR[15]  (.D(test_0_HADDR[15]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[15]));
    SLE \regHADDR[10]  (.D(test_0_HADDR[10]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[10]));
    SLE \regHADDR[6]  (.D(test_0_HADDR[6]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[6]));
    SLE \regHADDR[9]  (.D(test_0_HADDR[9]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[9]));
    SLE \regHADDR[8]  (.D(test_0_HADDR[8]), .CLK(GL0_INST), .EN(
        masterAddrClockEnable_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(regHADDR[8]));
    
endmodule


module COREAHBLITE_SLAVEARBITER_Z3_1(
       masterAddrInProg_0,
       M0GATEDHSIZE_0,
       N_128_i,
       CoreAHBLite_0_AHBmslave16_HREADY,
       m0s16AddrSel,
       d_masterRegAddrSel,
       VCC_0,
       VCC_0_reto,
       GL0_INST,
       u8_sb_0_HPMS_READY
    );
output masterAddrInProg_0;
input  M0GATEDHSIZE_0;
output N_128_i;
input  CoreAHBLite_0_AHBmslave16_HREADY;
input  m0s16AddrSel;
input  d_masterRegAddrSel;
input  VCC_0;
output VCC_0_reto;
input  GL0_INST;
input  u8_sb_0_HPMS_READY;

    wire \arbRegSMCurrentState[14]_net_1 , VCC_net_1, N_141_i, 
        GND_net_1, N_127_sn, N_143_i, \arbRegSMCurrentState[0]_net_1 , 
        N_119_i, \arbRegSMCurrentState[1]_net_1 , N_121_i, 
        \arbRegSMCurrentState[3]_net_1 , N_125_i, 
        \arbRegSMCurrentState[5]_net_1 , \arbRegSMCurrentStateoi[5] , 
        \arbRegSMCurrentState[6]_net_1 , N_129_i, N_125_sn, N_131_i, 
        \arbRegSMCurrentState[9]_net_1 , \arbRegSMCurrentStateoi[9] , 
        \arbRegSMCurrentState[10]_net_1 , N_135_i, N_126_sn, N_137_i, 
        \arbRegSMCurrentState[13]_net_1 , \arbRegSMCurrentStateoi[13] , 
        d_masterRegAddrSel_reto, N_123_i_reto, N_123_i, N_189, N_189oi, 
        MASTERADDRINPROG_N_4, N_153, N_159, N_164, N_152, 
        \arbRegSMCurrentState_ns_i_0[1]_net_1 , N_166, 
        \arbRegSMCurrentState_ns_i_1[1]_net_1 , 
        arbRegSMCurrentState_ret_4_RNO_0_net_1;
    
    SLE arbRegSMCurrentState_ret_4 (.D(N_123_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(N_123_i_reto));
    CFG4 #( .INIT(16'h0F0B) )  
        \arbRegSMCurrentState_ns_i_1_RNI7CLF[1]  (.A(N_123_i_reto), .B(
        N_153), .C(\arbRegSMCurrentState_ns_i_1[1]_net_1 ), .D(
        CoreAHBLite_0_AHBmslave16_HREADY), .Y(N_121_i));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[11]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_126_sn), .Y(N_137_i));
    SLE arbRegSMCurrentState_ret_2 (.D(VCC_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(VCC_0_reto));
    SLE \arbRegSMCurrentState[3]  (.D(N_125_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[3]_net_1 ));
    CFG3 #( .INIT(8'hAE) )  \arbRegSMCurrentState_ns[13]  (.A(
        \arbRegSMCurrentState[14]_net_1 ), .B(
        \arbRegSMCurrentState[13]_net_1 ), .C(m0s16AddrSel), .Y(
        \arbRegSMCurrentStateoi[13] ));
    CFG3 #( .INIT(8'hAE) )  \arbRegSMCurrentState_ns[9]  (.A(
        \arbRegSMCurrentState[10]_net_1 ), .B(
        \arbRegSMCurrentState[9]_net_1 ), .C(m0s16AddrSel), .Y(
        \arbRegSMCurrentStateoi[9] ));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[7]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_125_sn), .Y(N_131_i));
    SLE \arbRegSMCurrentState[10]  (.D(N_135_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[10]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hB) )  \arbRegSMCurrentState_ns_i_o2[1]  (.A(
        m0s16AddrSel), .B(\arbRegSMCurrentState[1]_net_1 ), .Y(N_153));
    CFG4 #( .INIT(16'h0C0D) )  \arbRegSMCurrentState_RNO[0]  (.A(
        M0GATEDHSIZE_0), .B(\arbRegSMCurrentState[0]_net_1 ), .C(
        CoreAHBLite_0_AHBmslave16_HREADY), .D(N_152), .Y(N_119_i));
    SLE \arbRegSMCurrentState[0]  (.D(N_119_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[0]_net_1 ));
    SLE \arbRegSMCurrentState[7]  (.D(N_131_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(N_125_sn));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[15]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_127_sn), .Y(N_143_i));
    SLE \arbRegSMCurrentState[14]  (.D(N_141_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[14]_net_1 ));
    SLE \arbRegSMCurrentState[6]  (.D(N_129_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[6]_net_1 ));
    CFG4 #( .INIT(16'hFF02) )  \arbRegSMCurrentState_ns_i_0[1]  (.A(
        N_189), .B(\arbRegSMCurrentState[0]_net_1 ), .C(N_123_i_reto), 
        .D(N_164), .Y(\arbRegSMCurrentState_ns_i_0[1]_net_1 ));
    SLE \arbRegSMCurrentState[1]  (.D(N_121_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \arbRegSMCurrentState_RNO[6]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_125_sn), .Y(N_129_i));
    CFG2 #( .INIT(4'h8) )  \arbRegSMCurrentState_RNO[10]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_126_sn), .Y(N_135_i));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hDF02) )  MASTERADDRINPROG_m5_0_m3 (.A(
        d_masterRegAddrSel_reto), .B(VCC_0_reto), .C(N_189), .D(
        N_123_i_reto), .Y(MASTERADDRINPROG_N_4));
    CFG4 #( .INIT(16'hFEEE) )  MASTERADDRINPROG_m5_0 (.A(
        \arbRegSMCurrentState[3]_net_1 ), .B(
        \arbRegSMCurrentState[0]_net_1 ), .C(MASTERADDRINPROG_N_4), .D(
        m0s16AddrSel), .Y(masterAddrInProg_0));
    CFG4 #( .INIT(16'h2031) )  arbRegSMCurrentState_ret_4_RNO_0 (.A(
        m0s16AddrSel), .B(CoreAHBLite_0_AHBmslave16_HREADY), .C(N_189), 
        .D(N_123_i_reto), .Y(arbRegSMCurrentState_ret_4_RNO_0_net_1));
    CFG2 #( .INIT(4'h8) )  \arbRegSMCurrentState_RNO[14]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_127_sn), .Y(N_141_i));
    SLE \arbRegSMCurrentState[9]  (.D(\arbRegSMCurrentStateoi[9] ), 
        .CLK(GL0_INST), .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\arbRegSMCurrentState[9]_net_1 ));
    CFG4 #( .INIT(16'hF2F0) )  \arbRegSMCurrentState_ns_i_1[1]  (.A(
        M0GATEDHSIZE_0), .B(\arbRegSMCurrentState[0]_net_1 ), .C(
        \arbRegSMCurrentState_ns_i_0[1]_net_1 ), .D(N_153), .Y(
        \arbRegSMCurrentState_ns_i_1[1]_net_1 ));
    SLE \arbRegSMCurrentState[13]  (.D(\arbRegSMCurrentStateoi[13] ), 
        .CLK(GL0_INST), .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\arbRegSMCurrentState[13]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \arbRegSMCurrentState_ns_i_a2_1[1]  (.A(
        \arbRegSMCurrentState[1]_net_1 ), .B(
        \arbRegSMCurrentState[0]_net_1 ), .C(N_123_i_reto), .D(
        m0s16AddrSel), .Y(N_164));
    SLE \arbRegSMCurrentState[11]  (.D(N_137_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(N_126_sn));
    CFG4 #( .INIT(16'hFFFE) )  \arbRegSMCurrentState_RNIEHSU[7]  (.A(
        N_127_sn), .B(N_126_sn), .C(N_125_sn), .D(masterAddrInProg_0), 
        .Y(N_128_i));
    CFG4 #( .INIT(16'h0001) )  \arbRegSMCurrentState_ns_i_a2_3[1]  (.A(
        \arbRegSMCurrentStateoi[13] ), .B(\arbRegSMCurrentStateoi[9] ), 
        .C(\arbRegSMCurrentStateoi[5] ), .D(N_121_i), .Y(N_189oi));
    CFG2 #( .INIT(4'h7) )  \arbRegSMCurrentState_ns_i_o2[3]  (.A(
        m0s16AddrSel), .B(M0GATEDHSIZE_0), .Y(N_159));
    CFG2 #( .INIT(4'hD) )  \arbRegSMCurrentState_ns_i_o2[0]  (.A(
        m0s16AddrSel), .B(N_189), .Y(N_152));
    SLE \arbRegSMCurrentState[5]  (.D(\arbRegSMCurrentStateoi[5] ), 
        .CLK(GL0_INST), .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\arbRegSMCurrentState[5]_net_1 ));
    SLE \arbRegSMCurrentState[15]  (.D(N_143_i), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(N_127_sn));
    CFG3 #( .INIT(8'h02) )  \arbRegSMCurrentState_ns_i_a2[2]  (.A(
        N_152), .B(\arbRegSMCurrentState[3]_net_1 ), .C(N_123_i_reto), 
        .Y(N_166));
    SLE arbRegSMCurrentState_ret_5 (.D(N_189oi), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(N_189));
    CFG3 #( .INIT(8'hAE) )  \arbRegSMCurrentState_ns[5]  (.A(
        \arbRegSMCurrentState[6]_net_1 ), .B(
        \arbRegSMCurrentState[5]_net_1 ), .C(m0s16AddrSel), .Y(
        \arbRegSMCurrentStateoi[5] ));
    CFG4 #( .INIT(16'h000E) )  arbRegSMCurrentState_ret_4_RNO (.A(
        \arbRegSMCurrentState[3]_net_1 ), .B(M0GATEDHSIZE_0), .C(N_166)
        , .D(arbRegSMCurrentState_ret_4_RNO_0_net_1), .Y(N_123_i));
    SLE arbRegSMCurrentState_ret_3 (.D(d_masterRegAddrSel), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(d_masterRegAddrSel_reto));
    CFG4 #( .INIT(16'h0C0E) )  \arbRegSMCurrentState_RNO[3]  (.A(
        N_123_i_reto), .B(\arbRegSMCurrentState[3]_net_1 ), .C(
        CoreAHBLite_0_AHBmslave16_HREADY), .D(N_159), .Y(N_125_i));
    
endmodule


module COREAHBLITE_SLAVESTAGE_0s_0_0_0(
       regHADDR,
       test_0_HADDR,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       test_0_HWDATA,
       CoreAHBLite_0_AHBmslave16_HADDR_28,
       CoreAHBLite_0_AHBmslave16_HADDR_27,
       CoreAHBLite_0_AHBmslave16_HADDR_14,
       CoreAHBLite_0_AHBmslave16_HADDR_0,
       CoreAHBLite_0_AHBmslave16_HADDR_1,
       CoreAHBLite_0_AHBmslave16_HADDR_2,
       CoreAHBLite_0_AHBmslave16_HADDR_3,
       CoreAHBLite_0_AHBmslave16_HADDR_4,
       CoreAHBLite_0_AHBmslave16_HADDR_5,
       CoreAHBLite_0_AHBmslave16_HADDR_6,
       CoreAHBLite_0_AHBmslave16_HADDR_7,
       CoreAHBLite_0_AHBmslave16_HADDR_8,
       CoreAHBLite_0_AHBmslave16_HADDR_9,
       CoreAHBLite_0_AHBmslave16_HADDR_10,
       CoreAHBLite_0_AHBmslave16_HADDR_11,
       CoreAHBLite_0_AHBmslave16_HADDR_12,
       CoreAHBLite_0_AHBmslave16_HADDR_13,
       CoreAHBLite_0_AHBmslave16_HTRANS_0,
       CoreAHBLite_0_AHBmslave16_HSIZE_0,
       M0GATEDHSIZE_0,
       M0GATEDHADDR_0,
       M0GATEDHADDR_13,
       masterAddrInProg_0,
       masterDataInProg_0,
       VCC_0_reto,
       VCC_0,
       d_masterRegAddrSel,
       N_128_i,
       CoreAHBLite_0_AHBmslave16_HWRITE,
       masterRegAddrSel,
       regHWRITE,
       test_0_HWRITE,
       m0s16AddrSel,
       CoreAHBLite_0_AHBmslave16_HREADY,
       GL0_INST,
       u8_sb_0_HPMS_READY
    );
input  [15:2] regHADDR;
input  [15:2] test_0_HADDR;
output [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
input  [31:0] test_0_HWDATA;
output CoreAHBLite_0_AHBmslave16_HADDR_28;
output CoreAHBLite_0_AHBmslave16_HADDR_27;
output CoreAHBLite_0_AHBmslave16_HADDR_14;
output CoreAHBLite_0_AHBmslave16_HADDR_0;
output CoreAHBLite_0_AHBmslave16_HADDR_1;
output CoreAHBLite_0_AHBmslave16_HADDR_2;
output CoreAHBLite_0_AHBmslave16_HADDR_3;
output CoreAHBLite_0_AHBmslave16_HADDR_4;
output CoreAHBLite_0_AHBmslave16_HADDR_5;
output CoreAHBLite_0_AHBmslave16_HADDR_6;
output CoreAHBLite_0_AHBmslave16_HADDR_7;
output CoreAHBLite_0_AHBmslave16_HADDR_8;
output CoreAHBLite_0_AHBmslave16_HADDR_9;
output CoreAHBLite_0_AHBmslave16_HADDR_10;
output CoreAHBLite_0_AHBmslave16_HADDR_11;
output CoreAHBLite_0_AHBmslave16_HADDR_12;
output CoreAHBLite_0_AHBmslave16_HADDR_13;
output CoreAHBLite_0_AHBmslave16_HTRANS_0;
output CoreAHBLite_0_AHBmslave16_HSIZE_0;
input  M0GATEDHSIZE_0;
input  M0GATEDHADDR_0;
input  M0GATEDHADDR_13;
output masterAddrInProg_0;
output masterDataInProg_0;
output VCC_0_reto;
input  VCC_0;
input  d_masterRegAddrSel;
output N_128_i;
output CoreAHBLite_0_AHBmslave16_HWRITE;
input  masterRegAddrSel;
input  regHWRITE;
input  test_0_HWRITE;
input  m0s16AddrSel;
input  CoreAHBLite_0_AHBmslave16_HREADY;
input  GL0_INST;
input  u8_sb_0_HPMS_READY;

    wire VCC_net_1, masterDataInProg_55_net_1, GND_net_1;
    
    CFG4 #( .INIT(16'hCA00) )  HWRITE (.A(test_0_HWRITE), .B(regHWRITE)
        , .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HWRITE));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[4]  (.A(test_0_HADDR[4]), .B(
        regHADDR[4]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_2));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[5]  (.A(test_0_HADDR[5]), .B(
        regHADDR[5]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_3));
    CFG2 #( .INIT(4'h8) )  \HADDR[30]  (.A(masterAddrInProg_0), .B(
        M0GATEDHADDR_0), .Y(CoreAHBLite_0_AHBmslave16_HADDR_28));
    CFG2 #( .INIT(4'h8) )  \HWDATA[22]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[22]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[22]));
    CFG2 #( .INIT(4'h8) )  HTRANS (.A(masterAddrInProg_0), .B(
        m0s16AddrSel), .Y(CoreAHBLite_0_AHBmslave16_HTRANS_0));
    CFG2 #( .INIT(4'h8) )  \HWDATA[20]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[20]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[20]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[23]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[23]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[23]));
    CFG2 #( .INIT(4'h8) )  HMASTLOCK (.A(masterAddrInProg_0), .B(
        M0GATEDHSIZE_0), .Y(CoreAHBLite_0_AHBmslave16_HSIZE_0));
    CFG2 #( .INIT(4'h8) )  \HWDATA[12]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[12]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[12]));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  \HWDATA[29]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[29]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[29]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[10]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[10]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[10]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[31]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[31]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[31]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[13]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[13]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[13]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[10]  (.A(test_0_HADDR[10]), .B(
        regHADDR[10]), .C(masterRegAddrSel), .D(masterAddrInProg_0), 
        .Y(CoreAHBLite_0_AHBmslave16_HADDR_8));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[14]  (.A(test_0_HADDR[14]), .B(
        regHADDR[14]), .C(masterRegAddrSel), .D(masterAddrInProg_0), 
        .Y(CoreAHBLite_0_AHBmslave16_HADDR_12));
    CFG2 #( .INIT(4'h8) )  \HWDATA[0]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[0]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[0]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[4]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[4]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[4]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[28]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[28]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[28]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[19]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[19]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[19]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[15]  (.A(test_0_HADDR[15]), .B(
        regHADDR[15]), .C(masterRegAddrSel), .D(masterAddrInProg_0), 
        .Y(CoreAHBLite_0_AHBmslave16_HADDR_13));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[11]  (.A(test_0_HADDR[11]), .B(
        regHADDR[11]), .C(masterRegAddrSel), .D(masterAddrInProg_0), 
        .Y(CoreAHBLite_0_AHBmslave16_HADDR_9));
    CFG2 #( .INIT(4'h8) )  \HWDATA[25]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[25]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[25]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[24]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[24]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[24]));
    CFG2 #( .INIT(4'h8) )  \HADDR[16]  (.A(masterAddrInProg_0), .B(
        M0GATEDHADDR_0), .Y(CoreAHBLite_0_AHBmslave16_HADDR_14));
    CFG2 #( .INIT(4'h8) )  \HWDATA[27]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[27]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[27]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[18]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[18]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[18]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[3]  (.A(test_0_HADDR[3]), .B(
        regHADDR[3]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_1));
    GND GND (.Y(GND_net_1));
    SLE \masterDataInProg[0]  (.D(masterDataInProg_55_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(masterDataInProg_0));
    CFG2 #( .INIT(4'h8) )  \HWDATA[15]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[15]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[15]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[14]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[14]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[14]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[8]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[8]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[8]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[6]  (.A(test_0_HADDR[6]), .B(
        regHADDR[6]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_4));
    CFG2 #( .INIT(4'h8) )  \HWDATA[3]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[3]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[3]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[17]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[17]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[17]));
    CFG2 #( .INIT(4'h8) )  \HADDR[29]  (.A(masterAddrInProg_0), .B(
        M0GATEDHADDR_13), .Y(CoreAHBLite_0_AHBmslave16_HADDR_27));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[7]  (.A(test_0_HADDR[7]), .B(
        regHADDR[7]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_5));
    CFG2 #( .INIT(4'h8) )  \HWDATA[5]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[5]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[5]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[12]  (.A(test_0_HADDR[12]), .B(
        regHADDR[12]), .C(masterRegAddrSel), .D(masterAddrInProg_0), 
        .Y(CoreAHBLite_0_AHBmslave16_HADDR_10));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[13]  (.A(test_0_HADDR[13]), .B(
        regHADDR[13]), .C(masterRegAddrSel), .D(masterAddrInProg_0), 
        .Y(CoreAHBLite_0_AHBmslave16_HADDR_11));
    CFG3 #( .INIT(8'hB8) )  masterDataInProg_55 (.A(masterAddrInProg_0)
        , .B(CoreAHBLite_0_AHBmslave16_HREADY), .C(masterDataInProg_0), 
        .Y(masterDataInProg_55_net_1));
    CFG2 #( .INIT(4'h8) )  \HWDATA[30]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[30]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[30]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[9]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[9]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[9]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[7]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[7]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[7]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[1]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[1]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[1]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[6]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[6]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[6]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[8]  (.A(test_0_HADDR[8]), .B(
        regHADDR[8]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_6));
    COREAHBLITE_SLAVEARBITER_Z3_1 slave_arbiter (.masterAddrInProg_0(
        masterAddrInProg_0), .M0GATEDHSIZE_0(M0GATEDHSIZE_0), .N_128_i(
        N_128_i), .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .m0s16AddrSel(m0s16AddrSel), 
        .d_masterRegAddrSel(d_masterRegAddrSel), .VCC_0(VCC_0), 
        .VCC_0_reto(VCC_0_reto), .GL0_INST(GL0_INST), 
        .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY));
    CFG2 #( .INIT(4'h8) )  \HWDATA[21]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[21]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[21]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[26]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[26]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[26]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[9]  (.A(test_0_HADDR[9]), .B(
        regHADDR[9]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_7));
    CFG2 #( .INIT(4'h8) )  \HWDATA[2]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[2]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[2]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[11]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[11]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[11]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[16]  (.A(masterDataInProg_0), .B(
        test_0_HWDATA[16]), .Y(CoreAHBLite_0_AHBmslave16_HWDATA[16]));
    CFG4 #( .INIT(16'hCA00) )  \HADDR[2]  (.A(test_0_HADDR[2]), .B(
        regHADDR[2]), .C(masterRegAddrSel), .D(masterAddrInProg_0), .Y(
        CoreAHBLite_0_AHBmslave16_HADDR_0));
    
endmodule


module COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0_0s(
       test_0_HWDATA,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       test_0_HADDR,
       masterAddrInProg_0,
       CoreAHBLite_0_AHBmslave16_HSIZE_0,
       CoreAHBLite_0_AHBmslave16_HTRANS_0,
       CoreAHBLite_0_AHBmslave16_HADDR_28,
       CoreAHBLite_0_AHBmslave16_HADDR_27,
       CoreAHBLite_0_AHBmslave16_HADDR_14,
       CoreAHBLite_0_AHBmslave16_HADDR_0,
       CoreAHBLite_0_AHBmslave16_HADDR_1,
       CoreAHBLite_0_AHBmslave16_HADDR_2,
       CoreAHBLite_0_AHBmslave16_HADDR_3,
       CoreAHBLite_0_AHBmslave16_HADDR_4,
       CoreAHBLite_0_AHBmslave16_HADDR_5,
       CoreAHBLite_0_AHBmslave16_HADDR_6,
       CoreAHBLite_0_AHBmslave16_HADDR_7,
       CoreAHBLite_0_AHBmslave16_HADDR_8,
       CoreAHBLite_0_AHBmslave16_HADDR_9,
       CoreAHBLite_0_AHBmslave16_HADDR_10,
       CoreAHBLite_0_AHBmslave16_HADDR_11,
       CoreAHBLite_0_AHBmslave16_HADDR_12,
       CoreAHBLite_0_AHBmslave16_HADDR_13,
       test_0_HADDR_i_0,
       test_0_HTRANS_0,
       CoreAHBLite_0_AHBmslave16_HWRITE,
       N_128_i,
       u8_sb_0_HPMS_READY,
       GL0_INST,
       m0s16DataSel,
       test_0_HWRITE,
       CoreAHBLite_0_AHBmslave16_HREADY,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       CoreAHBLite_0_AHBmslave16_HREADY_m_0
    );
input  [31:0] test_0_HWDATA;
output [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
input  [16:2] test_0_HADDR;
output masterAddrInProg_0;
output CoreAHBLite_0_AHBmslave16_HSIZE_0;
output CoreAHBLite_0_AHBmslave16_HTRANS_0;
output CoreAHBLite_0_AHBmslave16_HADDR_28;
output CoreAHBLite_0_AHBmslave16_HADDR_27;
output CoreAHBLite_0_AHBmslave16_HADDR_14;
output CoreAHBLite_0_AHBmslave16_HADDR_0;
output CoreAHBLite_0_AHBmslave16_HADDR_1;
output CoreAHBLite_0_AHBmslave16_HADDR_2;
output CoreAHBLite_0_AHBmslave16_HADDR_3;
output CoreAHBLite_0_AHBmslave16_HADDR_4;
output CoreAHBLite_0_AHBmslave16_HADDR_5;
output CoreAHBLite_0_AHBmslave16_HADDR_6;
output CoreAHBLite_0_AHBmslave16_HADDR_7;
output CoreAHBLite_0_AHBmslave16_HADDR_8;
output CoreAHBLite_0_AHBmslave16_HADDR_9;
output CoreAHBLite_0_AHBmslave16_HADDR_10;
output CoreAHBLite_0_AHBmslave16_HADDR_11;
output CoreAHBLite_0_AHBmslave16_HADDR_12;
output CoreAHBLite_0_AHBmslave16_HADDR_13;
input  test_0_HADDR_i_0;
input  test_0_HTRANS_0;
output CoreAHBLite_0_AHBmslave16_HWRITE;
output N_128_i;
input  u8_sb_0_HPMS_READY;
input  GL0_INST;
output m0s16DataSel;
input  test_0_HWRITE;
input  CoreAHBLite_0_AHBmslave16_HREADY;
output u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
input  CoreAHBLite_0_AHBmslave16_HREADY_m_0;

    wire \masterDataInProg[0] , \M0GATEDHADDR[16] , \M0GATEDHADDR[29] , 
        \M0GATEDHSIZE[1] , \regHADDR[2] , \regHADDR[3] , \regHADDR[4] , 
        \regHADDR[5] , \regHADDR[6] , \regHADDR[7] , \regHADDR[8] , 
        \regHADDR[9] , \regHADDR[10] , \regHADDR[11] , \regHADDR[12] , 
        \regHADDR[13] , \regHADDR[14] , \regHADDR[15] , m0s16AddrSel, 
        VCC_0, VCC_0_reto, d_masterRegAddrSel, masterRegAddrSel, 
        regHWRITE, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    COREAHBLITE_MASTERSTAGE_1_1_85_65536_0s_0_1_0 masterstage_0 (
        .test_0_HADDR({test_0_HADDR[16], test_0_HADDR[15], 
        test_0_HADDR[14], test_0_HADDR[13], test_0_HADDR[12], 
        test_0_HADDR[11], test_0_HADDR[10], test_0_HADDR[9], 
        test_0_HADDR[8], test_0_HADDR[7], test_0_HADDR[6], 
        test_0_HADDR[5], test_0_HADDR[4], test_0_HADDR[3], 
        test_0_HADDR[2]}), .regHADDR({\regHADDR[15] , \regHADDR[14] , 
        \regHADDR[13] , \regHADDR[12] , \regHADDR[11] , \regHADDR[10] , 
        \regHADDR[9] , \regHADDR[8] , \regHADDR[7] , \regHADDR[6] , 
        \regHADDR[5] , \regHADDR[4] , \regHADDR[3] , \regHADDR[2] }), 
        .masterDataInProg_0(\masterDataInProg[0] ), .M0GATEDHADDR_0(
        \M0GATEDHADDR[16] ), .M0GATEDHADDR_13(\M0GATEDHADDR[29] ), 
        .test_0_HTRANS_0(test_0_HTRANS_0), .M0GATEDHSIZE_0(
        \M0GATEDHSIZE[1] ), .test_0_HADDR_i_0(test_0_HADDR_i_0), 
        .CoreAHBLite_0_AHBmslave16_HREADY_m_0(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .m0s16AddrSel(m0s16AddrSel), 
        .VCC_0(VCC_0), .VCC_0_reto(VCC_0_reto), .d_masterRegAddrSel(
        d_masterRegAddrSel), .masterRegAddrSel(masterRegAddrSel), 
        .test_0_HWRITE(test_0_HWRITE), .regHWRITE(regHWRITE), 
        .m0s16DataSel(m0s16DataSel), .GL0_INST(GL0_INST), 
        .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY));
    COREAHBLITE_SLAVESTAGE_0s_0_0_0 slavestage_16 (.regHADDR({
        \regHADDR[15] , \regHADDR[14] , \regHADDR[13] , \regHADDR[12] , 
        \regHADDR[11] , \regHADDR[10] , \regHADDR[9] , \regHADDR[8] , 
        \regHADDR[7] , \regHADDR[6] , \regHADDR[5] , \regHADDR[4] , 
        \regHADDR[3] , \regHADDR[2] }), .test_0_HADDR({
        test_0_HADDR[15], test_0_HADDR[14], test_0_HADDR[13], 
        test_0_HADDR[12], test_0_HADDR[11], test_0_HADDR[10], 
        test_0_HADDR[9], test_0_HADDR[8], test_0_HADDR[7], 
        test_0_HADDR[6], test_0_HADDR[5], test_0_HADDR[4], 
        test_0_HADDR[3], test_0_HADDR[2]}), 
        .CoreAHBLite_0_AHBmslave16_HWDATA({
        CoreAHBLite_0_AHBmslave16_HWDATA[31], 
        CoreAHBLite_0_AHBmslave16_HWDATA[30], 
        CoreAHBLite_0_AHBmslave16_HWDATA[29], 
        CoreAHBLite_0_AHBmslave16_HWDATA[28], 
        CoreAHBLite_0_AHBmslave16_HWDATA[27], 
        CoreAHBLite_0_AHBmslave16_HWDATA[26], 
        CoreAHBLite_0_AHBmslave16_HWDATA[25], 
        CoreAHBLite_0_AHBmslave16_HWDATA[24], 
        CoreAHBLite_0_AHBmslave16_HWDATA[23], 
        CoreAHBLite_0_AHBmslave16_HWDATA[22], 
        CoreAHBLite_0_AHBmslave16_HWDATA[21], 
        CoreAHBLite_0_AHBmslave16_HWDATA[20], 
        CoreAHBLite_0_AHBmslave16_HWDATA[19], 
        CoreAHBLite_0_AHBmslave16_HWDATA[18], 
        CoreAHBLite_0_AHBmslave16_HWDATA[17], 
        CoreAHBLite_0_AHBmslave16_HWDATA[16], 
        CoreAHBLite_0_AHBmslave16_HWDATA[15], 
        CoreAHBLite_0_AHBmslave16_HWDATA[14], 
        CoreAHBLite_0_AHBmslave16_HWDATA[13], 
        CoreAHBLite_0_AHBmslave16_HWDATA[12], 
        CoreAHBLite_0_AHBmslave16_HWDATA[11], 
        CoreAHBLite_0_AHBmslave16_HWDATA[10], 
        CoreAHBLite_0_AHBmslave16_HWDATA[9], 
        CoreAHBLite_0_AHBmslave16_HWDATA[8], 
        CoreAHBLite_0_AHBmslave16_HWDATA[7], 
        CoreAHBLite_0_AHBmslave16_HWDATA[6], 
        CoreAHBLite_0_AHBmslave16_HWDATA[5], 
        CoreAHBLite_0_AHBmslave16_HWDATA[4], 
        CoreAHBLite_0_AHBmslave16_HWDATA[3], 
        CoreAHBLite_0_AHBmslave16_HWDATA[2], 
        CoreAHBLite_0_AHBmslave16_HWDATA[1], 
        CoreAHBLite_0_AHBmslave16_HWDATA[0]}), .test_0_HWDATA({
        test_0_HWDATA[31], test_0_HWDATA[30], test_0_HWDATA[29], 
        test_0_HWDATA[28], test_0_HWDATA[27], test_0_HWDATA[26], 
        test_0_HWDATA[25], test_0_HWDATA[24], test_0_HWDATA[23], 
        test_0_HWDATA[22], test_0_HWDATA[21], test_0_HWDATA[20], 
        test_0_HWDATA[19], test_0_HWDATA[18], test_0_HWDATA[17], 
        test_0_HWDATA[16], test_0_HWDATA[15], test_0_HWDATA[14], 
        test_0_HWDATA[13], test_0_HWDATA[12], test_0_HWDATA[11], 
        test_0_HWDATA[10], test_0_HWDATA[9], test_0_HWDATA[8], 
        test_0_HWDATA[7], test_0_HWDATA[6], test_0_HWDATA[5], 
        test_0_HWDATA[4], test_0_HWDATA[3], test_0_HWDATA[2], 
        test_0_HWDATA[1], test_0_HWDATA[0]}), 
        .CoreAHBLite_0_AHBmslave16_HADDR_28(
        CoreAHBLite_0_AHBmslave16_HADDR_28), 
        .CoreAHBLite_0_AHBmslave16_HADDR_27(
        CoreAHBLite_0_AHBmslave16_HADDR_27), 
        .CoreAHBLite_0_AHBmslave16_HADDR_14(
        CoreAHBLite_0_AHBmslave16_HADDR_14), 
        .CoreAHBLite_0_AHBmslave16_HADDR_0(
        CoreAHBLite_0_AHBmslave16_HADDR_0), 
        .CoreAHBLite_0_AHBmslave16_HADDR_1(
        CoreAHBLite_0_AHBmslave16_HADDR_1), 
        .CoreAHBLite_0_AHBmslave16_HADDR_2(
        CoreAHBLite_0_AHBmslave16_HADDR_2), 
        .CoreAHBLite_0_AHBmslave16_HADDR_3(
        CoreAHBLite_0_AHBmslave16_HADDR_3), 
        .CoreAHBLite_0_AHBmslave16_HADDR_4(
        CoreAHBLite_0_AHBmslave16_HADDR_4), 
        .CoreAHBLite_0_AHBmslave16_HADDR_5(
        CoreAHBLite_0_AHBmslave16_HADDR_5), 
        .CoreAHBLite_0_AHBmslave16_HADDR_6(
        CoreAHBLite_0_AHBmslave16_HADDR_6), 
        .CoreAHBLite_0_AHBmslave16_HADDR_7(
        CoreAHBLite_0_AHBmslave16_HADDR_7), 
        .CoreAHBLite_0_AHBmslave16_HADDR_8(
        CoreAHBLite_0_AHBmslave16_HADDR_8), 
        .CoreAHBLite_0_AHBmslave16_HADDR_9(
        CoreAHBLite_0_AHBmslave16_HADDR_9), 
        .CoreAHBLite_0_AHBmslave16_HADDR_10(
        CoreAHBLite_0_AHBmslave16_HADDR_10), 
        .CoreAHBLite_0_AHBmslave16_HADDR_11(
        CoreAHBLite_0_AHBmslave16_HADDR_11), 
        .CoreAHBLite_0_AHBmslave16_HADDR_12(
        CoreAHBLite_0_AHBmslave16_HADDR_12), 
        .CoreAHBLite_0_AHBmslave16_HADDR_13(
        CoreAHBLite_0_AHBmslave16_HADDR_13), 
        .CoreAHBLite_0_AHBmslave16_HTRANS_0(
        CoreAHBLite_0_AHBmslave16_HTRANS_0), 
        .CoreAHBLite_0_AHBmslave16_HSIZE_0(
        CoreAHBLite_0_AHBmslave16_HSIZE_0), .M0GATEDHSIZE_0(
        \M0GATEDHSIZE[1] ), .M0GATEDHADDR_0(\M0GATEDHADDR[16] ), 
        .M0GATEDHADDR_13(\M0GATEDHADDR[29] ), .masterAddrInProg_0(
        masterAddrInProg_0), .masterDataInProg_0(\masterDataInProg[0] )
        , .VCC_0_reto(VCC_0_reto), .VCC_0(VCC_0), .d_masterRegAddrSel(
        d_masterRegAddrSel), .N_128_i(N_128_i), 
        .CoreAHBLite_0_AHBmslave16_HWRITE(
        CoreAHBLite_0_AHBmslave16_HWRITE), .masterRegAddrSel(
        masterRegAddrSel), .regHWRITE(regHWRITE), .test_0_HWRITE(
        test_0_HWRITE), .m0s16AddrSel(m0s16AddrSel), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .GL0_INST(GL0_INST), 
        .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY));
    
endmodule


module CoreAHBLite_Z4(
       test_0_HADDR,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       test_0_HWDATA,
       test_0_HTRANS_0,
       test_0_HADDR_i_0,
       CoreAHBLite_0_AHBmslave16_HADDR_28,
       CoreAHBLite_0_AHBmslave16_HADDR_27,
       CoreAHBLite_0_AHBmslave16_HADDR_14,
       CoreAHBLite_0_AHBmslave16_HADDR_0,
       CoreAHBLite_0_AHBmslave16_HADDR_1,
       CoreAHBLite_0_AHBmslave16_HADDR_2,
       CoreAHBLite_0_AHBmslave16_HADDR_3,
       CoreAHBLite_0_AHBmslave16_HADDR_4,
       CoreAHBLite_0_AHBmslave16_HADDR_5,
       CoreAHBLite_0_AHBmslave16_HADDR_6,
       CoreAHBLite_0_AHBmslave16_HADDR_7,
       CoreAHBLite_0_AHBmslave16_HADDR_8,
       CoreAHBLite_0_AHBmslave16_HADDR_9,
       CoreAHBLite_0_AHBmslave16_HADDR_10,
       CoreAHBLite_0_AHBmslave16_HADDR_11,
       CoreAHBLite_0_AHBmslave16_HADDR_12,
       CoreAHBLite_0_AHBmslave16_HADDR_13,
       CoreAHBLite_0_AHBmslave16_HTRANS_0,
       CoreAHBLite_0_AHBmslave16_HSIZE_0,
       masterAddrInProg_0,
       CoreAHBLite_0_AHBmslave16_HREADY_m_0,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       CoreAHBLite_0_AHBmslave16_HREADY,
       test_0_HWRITE,
       m0s16DataSel,
       GL0_INST,
       u8_sb_0_HPMS_READY,
       N_128_i,
       CoreAHBLite_0_AHBmslave16_HWRITE
    );
input  [16:2] test_0_HADDR;
output [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
input  [31:0] test_0_HWDATA;
input  test_0_HTRANS_0;
input  test_0_HADDR_i_0;
output CoreAHBLite_0_AHBmslave16_HADDR_28;
output CoreAHBLite_0_AHBmslave16_HADDR_27;
output CoreAHBLite_0_AHBmslave16_HADDR_14;
output CoreAHBLite_0_AHBmslave16_HADDR_0;
output CoreAHBLite_0_AHBmslave16_HADDR_1;
output CoreAHBLite_0_AHBmslave16_HADDR_2;
output CoreAHBLite_0_AHBmslave16_HADDR_3;
output CoreAHBLite_0_AHBmslave16_HADDR_4;
output CoreAHBLite_0_AHBmslave16_HADDR_5;
output CoreAHBLite_0_AHBmslave16_HADDR_6;
output CoreAHBLite_0_AHBmslave16_HADDR_7;
output CoreAHBLite_0_AHBmslave16_HADDR_8;
output CoreAHBLite_0_AHBmslave16_HADDR_9;
output CoreAHBLite_0_AHBmslave16_HADDR_10;
output CoreAHBLite_0_AHBmslave16_HADDR_11;
output CoreAHBLite_0_AHBmslave16_HADDR_12;
output CoreAHBLite_0_AHBmslave16_HADDR_13;
output CoreAHBLite_0_AHBmslave16_HTRANS_0;
output CoreAHBLite_0_AHBmslave16_HSIZE_0;
output masterAddrInProg_0;
input  CoreAHBLite_0_AHBmslave16_HREADY_m_0;
output u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
input  CoreAHBLite_0_AHBmslave16_HREADY;
input  test_0_HWRITE;
output m0s16DataSel;
input  GL0_INST;
input  u8_sb_0_HPMS_READY;
output N_128_i;
output CoreAHBLite_0_AHBmslave16_HWRITE;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0_0s matrix4x16 (
        .test_0_HWDATA({test_0_HWDATA[31], test_0_HWDATA[30], 
        test_0_HWDATA[29], test_0_HWDATA[28], test_0_HWDATA[27], 
        test_0_HWDATA[26], test_0_HWDATA[25], test_0_HWDATA[24], 
        test_0_HWDATA[23], test_0_HWDATA[22], test_0_HWDATA[21], 
        test_0_HWDATA[20], test_0_HWDATA[19], test_0_HWDATA[18], 
        test_0_HWDATA[17], test_0_HWDATA[16], test_0_HWDATA[15], 
        test_0_HWDATA[14], test_0_HWDATA[13], test_0_HWDATA[12], 
        test_0_HWDATA[11], test_0_HWDATA[10], test_0_HWDATA[9], 
        test_0_HWDATA[8], test_0_HWDATA[7], test_0_HWDATA[6], 
        test_0_HWDATA[5], test_0_HWDATA[4], test_0_HWDATA[3], 
        test_0_HWDATA[2], test_0_HWDATA[1], test_0_HWDATA[0]}), 
        .CoreAHBLite_0_AHBmslave16_HWDATA({
        CoreAHBLite_0_AHBmslave16_HWDATA[31], 
        CoreAHBLite_0_AHBmslave16_HWDATA[30], 
        CoreAHBLite_0_AHBmslave16_HWDATA[29], 
        CoreAHBLite_0_AHBmslave16_HWDATA[28], 
        CoreAHBLite_0_AHBmslave16_HWDATA[27], 
        CoreAHBLite_0_AHBmslave16_HWDATA[26], 
        CoreAHBLite_0_AHBmslave16_HWDATA[25], 
        CoreAHBLite_0_AHBmslave16_HWDATA[24], 
        CoreAHBLite_0_AHBmslave16_HWDATA[23], 
        CoreAHBLite_0_AHBmslave16_HWDATA[22], 
        CoreAHBLite_0_AHBmslave16_HWDATA[21], 
        CoreAHBLite_0_AHBmslave16_HWDATA[20], 
        CoreAHBLite_0_AHBmslave16_HWDATA[19], 
        CoreAHBLite_0_AHBmslave16_HWDATA[18], 
        CoreAHBLite_0_AHBmslave16_HWDATA[17], 
        CoreAHBLite_0_AHBmslave16_HWDATA[16], 
        CoreAHBLite_0_AHBmslave16_HWDATA[15], 
        CoreAHBLite_0_AHBmslave16_HWDATA[14], 
        CoreAHBLite_0_AHBmslave16_HWDATA[13], 
        CoreAHBLite_0_AHBmslave16_HWDATA[12], 
        CoreAHBLite_0_AHBmslave16_HWDATA[11], 
        CoreAHBLite_0_AHBmslave16_HWDATA[10], 
        CoreAHBLite_0_AHBmslave16_HWDATA[9], 
        CoreAHBLite_0_AHBmslave16_HWDATA[8], 
        CoreAHBLite_0_AHBmslave16_HWDATA[7], 
        CoreAHBLite_0_AHBmslave16_HWDATA[6], 
        CoreAHBLite_0_AHBmslave16_HWDATA[5], 
        CoreAHBLite_0_AHBmslave16_HWDATA[4], 
        CoreAHBLite_0_AHBmslave16_HWDATA[3], 
        CoreAHBLite_0_AHBmslave16_HWDATA[2], 
        CoreAHBLite_0_AHBmslave16_HWDATA[1], 
        CoreAHBLite_0_AHBmslave16_HWDATA[0]}), .test_0_HADDR({
        test_0_HADDR[16], test_0_HADDR[15], test_0_HADDR[14], 
        test_0_HADDR[13], test_0_HADDR[12], test_0_HADDR[11], 
        test_0_HADDR[10], test_0_HADDR[9], test_0_HADDR[8], 
        test_0_HADDR[7], test_0_HADDR[6], test_0_HADDR[5], 
        test_0_HADDR[4], test_0_HADDR[3], test_0_HADDR[2]}), 
        .masterAddrInProg_0(masterAddrInProg_0), 
        .CoreAHBLite_0_AHBmslave16_HSIZE_0(
        CoreAHBLite_0_AHBmslave16_HSIZE_0), 
        .CoreAHBLite_0_AHBmslave16_HTRANS_0(
        CoreAHBLite_0_AHBmslave16_HTRANS_0), 
        .CoreAHBLite_0_AHBmslave16_HADDR_28(
        CoreAHBLite_0_AHBmslave16_HADDR_28), 
        .CoreAHBLite_0_AHBmslave16_HADDR_27(
        CoreAHBLite_0_AHBmslave16_HADDR_27), 
        .CoreAHBLite_0_AHBmslave16_HADDR_14(
        CoreAHBLite_0_AHBmslave16_HADDR_14), 
        .CoreAHBLite_0_AHBmslave16_HADDR_0(
        CoreAHBLite_0_AHBmslave16_HADDR_0), 
        .CoreAHBLite_0_AHBmslave16_HADDR_1(
        CoreAHBLite_0_AHBmslave16_HADDR_1), 
        .CoreAHBLite_0_AHBmslave16_HADDR_2(
        CoreAHBLite_0_AHBmslave16_HADDR_2), 
        .CoreAHBLite_0_AHBmslave16_HADDR_3(
        CoreAHBLite_0_AHBmslave16_HADDR_3), 
        .CoreAHBLite_0_AHBmslave16_HADDR_4(
        CoreAHBLite_0_AHBmslave16_HADDR_4), 
        .CoreAHBLite_0_AHBmslave16_HADDR_5(
        CoreAHBLite_0_AHBmslave16_HADDR_5), 
        .CoreAHBLite_0_AHBmslave16_HADDR_6(
        CoreAHBLite_0_AHBmslave16_HADDR_6), 
        .CoreAHBLite_0_AHBmslave16_HADDR_7(
        CoreAHBLite_0_AHBmslave16_HADDR_7), 
        .CoreAHBLite_0_AHBmslave16_HADDR_8(
        CoreAHBLite_0_AHBmslave16_HADDR_8), 
        .CoreAHBLite_0_AHBmslave16_HADDR_9(
        CoreAHBLite_0_AHBmslave16_HADDR_9), 
        .CoreAHBLite_0_AHBmslave16_HADDR_10(
        CoreAHBLite_0_AHBmslave16_HADDR_10), 
        .CoreAHBLite_0_AHBmslave16_HADDR_11(
        CoreAHBLite_0_AHBmslave16_HADDR_11), 
        .CoreAHBLite_0_AHBmslave16_HADDR_12(
        CoreAHBLite_0_AHBmslave16_HADDR_12), 
        .CoreAHBLite_0_AHBmslave16_HADDR_13(
        CoreAHBLite_0_AHBmslave16_HADDR_13), .test_0_HADDR_i_0(
        test_0_HADDR_i_0), .test_0_HTRANS_0(test_0_HTRANS_0), 
        .CoreAHBLite_0_AHBmslave16_HWRITE(
        CoreAHBLite_0_AHBmslave16_HWRITE), .N_128_i(N_128_i), 
        .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY), .GL0_INST(GL0_INST), 
        .m0s16DataSel(m0s16DataSel), .test_0_HWRITE(test_0_HWRITE), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), 
        .CoreAHBLite_0_AHBmslave16_HREADY_m_0(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0));
    GND GND (.Y(GND_net_1));
    
endmodule


module u8_sb_CCC_0_FCCC(
       u8_sb_0_FIC_0_LOCK,
       GL0_INST,
       mclk_c
    );
output u8_sb_0_FIC_0_LOCK;
output GL0_INST;
input  mclk_c;

    wire mclk_c_i, GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST_inst_1 (.A(GL0_net), .Y(GL0_INST));
    CFG1 #( .INIT(2'h1) )  CCC_INST_RNO (.A(mclk_c), .Y(mclk_c_i));
    CCC #( .INIT(210'h0000007FB8000045174000318C6318C1F18C61F00404040400101)
        , .VCOFREQUENCY(786.432) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(
        ), .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(
        u8_sb_0_FIC_0_LOCK), .BUSY(), .CLK0(mclk_c_i), .CLK1(VCC_net_1)
        , .CLK2(VCC_net_1), .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), 
        .NGMUX1_SEL(GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(
        GND_net_1), .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(
        VCC_net_1), .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(
        VCC_net_1), .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(
        VCC_net_1), .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(
        VCC_net_1), .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(GND_net_1), .RCOSC_1MHZ(GND_net_1), 
        .XTLOSC(GND_net_1));
    
endmodule


module u8_sb(
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0,
       test_0_HWDATA,
       test_0_HADDR,
       test_0_HADDR_i_0,
       test_0_HTRANS_0,
       u8_sb_0_HPMS_READY,
       test_0_HWRITE,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       mclk_c,
       DEVRST_N
    );
output [31:0] u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0;
input  [31:0] test_0_HWDATA;
input  [16:2] test_0_HADDR;
input  test_0_HADDR_i_0;
input  test_0_HTRANS_0;
output u8_sb_0_HPMS_READY;
input  test_0_HWRITE;
output u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
input  mclk_c;
input  DEVRST_N;

    wire SYSRESET_POR_net_1, u8_sb_0_FIC_0_LOCK, GL0_INST, 
        \CoreAHBLite_0_AHBmslave16_HADDR[30] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[29] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[16] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[2] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[3] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[4] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[5] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[6] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[7] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[8] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[9] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[10] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[11] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[12] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[13] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[14] , 
        \CoreAHBLite_0_AHBmslave16_HADDR[15] , 
        \CoreAHBLite_0_AHBmslave16_HTRANS[1] , 
        \CoreAHBLite_0_AHBmslave16_HSIZE[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[0] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[31] , \masterAddrInProg[0] , 
        CoreAHBLite_0_AHBmslave16_HREADY_m_0, 
        CoreAHBLite_0_AHBmslave16_HREADY, m0s16DataSel, N_128_i, 
        CoreAHBLite_0_AHBmslave16_HWRITE, 
        u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N, 
        u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F, GND_net_1, VCC_net_1;
    
    u8_sb_HPMS u8_sb_HPMS_0 (.CoreAHBLite_0_AHBmslave16_HWDATA({
        \CoreAHBLite_0_AHBmslave16_HWDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[0] }), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0({
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0]}), 
        .CoreAHBLite_0_AHBmslave16_HTRANS_0(
        \CoreAHBLite_0_AHBmslave16_HTRANS[1] ), 
        .CoreAHBLite_0_AHBmslave16_HSIZE_0(
        \CoreAHBLite_0_AHBmslave16_HSIZE[1] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_0(
        \CoreAHBLite_0_AHBmslave16_HADDR[2] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_1(
        \CoreAHBLite_0_AHBmslave16_HADDR[3] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_2(
        \CoreAHBLite_0_AHBmslave16_HADDR[4] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_3(
        \CoreAHBLite_0_AHBmslave16_HADDR[5] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_4(
        \CoreAHBLite_0_AHBmslave16_HADDR[6] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_5(
        \CoreAHBLite_0_AHBmslave16_HADDR[7] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_6(
        \CoreAHBLite_0_AHBmslave16_HADDR[8] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_7(
        \CoreAHBLite_0_AHBmslave16_HADDR[9] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_8(
        \CoreAHBLite_0_AHBmslave16_HADDR[10] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_9(
        \CoreAHBLite_0_AHBmslave16_HADDR[11] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_10(
        \CoreAHBLite_0_AHBmslave16_HADDR[12] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_11(
        \CoreAHBLite_0_AHBmslave16_HADDR[13] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_12(
        \CoreAHBLite_0_AHBmslave16_HADDR[14] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_13(
        \CoreAHBLite_0_AHBmslave16_HADDR[15] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_14(
        \CoreAHBLite_0_AHBmslave16_HADDR[16] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_27(
        \CoreAHBLite_0_AHBmslave16_HADDR[29] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_28(
        \CoreAHBLite_0_AHBmslave16_HADDR[30] ), .masterAddrInProg_0(
        \masterAddrInProg[0] ), .GL0_INST(GL0_INST), 
        .u8_sb_0_FIC_0_LOCK(u8_sb_0_FIC_0_LOCK), 
        .CoreAHBLite_0_AHBmslave16_HWRITE(
        CoreAHBLite_0_AHBmslave16_HWRITE), .N_128_i(N_128_i), 
        .u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F(
        u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F), 
        .u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N(
        u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), .m0s16DataSel(
        m0s16DataSel), .CoreAHBLite_0_AHBmslave16_HREADY_m_0(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY));
    CoreResetP_Z5 CORERESETP_0 (.u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N(
        u8_sb_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F(
        u8_sb_HPMS_TMP_0_MSS_RESET_N_M2F), .SYSRESET_POR(
        SYSRESET_POR_net_1), .GL0_INST(GL0_INST), .u8_sb_0_HPMS_READY(
        u8_sb_0_HPMS_READY));
    CoreAHBLite_Z4 CoreAHBLite_0 (.test_0_HADDR({test_0_HADDR[16], 
        test_0_HADDR[15], test_0_HADDR[14], test_0_HADDR[13], 
        test_0_HADDR[12], test_0_HADDR[11], test_0_HADDR[10], 
        test_0_HADDR[9], test_0_HADDR[8], test_0_HADDR[7], 
        test_0_HADDR[6], test_0_HADDR[5], test_0_HADDR[4], 
        test_0_HADDR[3], test_0_HADDR[2]}), 
        .CoreAHBLite_0_AHBmslave16_HWDATA({
        \CoreAHBLite_0_AHBmslave16_HWDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[0] }), .test_0_HWDATA({
        test_0_HWDATA[31], test_0_HWDATA[30], test_0_HWDATA[29], 
        test_0_HWDATA[28], test_0_HWDATA[27], test_0_HWDATA[26], 
        test_0_HWDATA[25], test_0_HWDATA[24], test_0_HWDATA[23], 
        test_0_HWDATA[22], test_0_HWDATA[21], test_0_HWDATA[20], 
        test_0_HWDATA[19], test_0_HWDATA[18], test_0_HWDATA[17], 
        test_0_HWDATA[16], test_0_HWDATA[15], test_0_HWDATA[14], 
        test_0_HWDATA[13], test_0_HWDATA[12], test_0_HWDATA[11], 
        test_0_HWDATA[10], test_0_HWDATA[9], test_0_HWDATA[8], 
        test_0_HWDATA[7], test_0_HWDATA[6], test_0_HWDATA[5], 
        test_0_HWDATA[4], test_0_HWDATA[3], test_0_HWDATA[2], 
        test_0_HWDATA[1], test_0_HWDATA[0]}), .test_0_HTRANS_0(
        test_0_HTRANS_0), .test_0_HADDR_i_0(test_0_HADDR_i_0), 
        .CoreAHBLite_0_AHBmslave16_HADDR_28(
        \CoreAHBLite_0_AHBmslave16_HADDR[30] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_27(
        \CoreAHBLite_0_AHBmslave16_HADDR[29] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_14(
        \CoreAHBLite_0_AHBmslave16_HADDR[16] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_0(
        \CoreAHBLite_0_AHBmslave16_HADDR[2] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_1(
        \CoreAHBLite_0_AHBmslave16_HADDR[3] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_2(
        \CoreAHBLite_0_AHBmslave16_HADDR[4] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_3(
        \CoreAHBLite_0_AHBmslave16_HADDR[5] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_4(
        \CoreAHBLite_0_AHBmslave16_HADDR[6] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_5(
        \CoreAHBLite_0_AHBmslave16_HADDR[7] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_6(
        \CoreAHBLite_0_AHBmslave16_HADDR[8] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_7(
        \CoreAHBLite_0_AHBmslave16_HADDR[9] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_8(
        \CoreAHBLite_0_AHBmslave16_HADDR[10] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_9(
        \CoreAHBLite_0_AHBmslave16_HADDR[11] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_10(
        \CoreAHBLite_0_AHBmslave16_HADDR[12] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_11(
        \CoreAHBLite_0_AHBmslave16_HADDR[13] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_12(
        \CoreAHBLite_0_AHBmslave16_HADDR[14] ), 
        .CoreAHBLite_0_AHBmslave16_HADDR_13(
        \CoreAHBLite_0_AHBmslave16_HADDR[15] ), 
        .CoreAHBLite_0_AHBmslave16_HTRANS_0(
        \CoreAHBLite_0_AHBmslave16_HTRANS[1] ), 
        .CoreAHBLite_0_AHBmslave16_HSIZE_0(
        \CoreAHBLite_0_AHBmslave16_HSIZE[1] ), .masterAddrInProg_0(
        \masterAddrInProg[0] ), .CoreAHBLite_0_AHBmslave16_HREADY_m_0(
        CoreAHBLite_0_AHBmslave16_HREADY_m_0), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .test_0_HWRITE(
        test_0_HWRITE), .m0s16DataSel(m0s16DataSel), .GL0_INST(
        GL0_INST), .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY), .N_128_i(
        N_128_i), .CoreAHBLite_0_AHBmslave16_HWRITE(
        CoreAHBLite_0_AHBmslave16_HWRITE));
    VCC VCC (.Y(VCC_net_1));
    u8_sb_CCC_0_FCCC CCC_0 (.u8_sb_0_FIC_0_LOCK(u8_sb_0_FIC_0_LOCK), 
        .GL0_INST(GL0_INST), .mclk_c(mclk_c));
    GND GND (.Y(GND_net_1));
    SYSRESET SYSRESET_POR (.POWER_ON_RESET_N(SYSRESET_POR_net_1), 
        .DEVRST_N(DEVRST_N));
    
endmodule


module crc7(
       crc,
       bit,
       crc_en,
       sdclk_n_1,
       crc_clr_i
    );
output [6:0] crc;
input  bit;
input  crc_en;
input  sdclk_n_1;
input  crc_clr_i;

    wire VCC_net_1, GND_net_1, N_110_i_i, N_94_i;
    
    SLE \CRC[6]  (.D(crc[5]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[6]));
    SLE \CRC[1]  (.D(crc[0]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[1]));
    CFG2 #( .INIT(4'h6) )  inv_0_x2 (.A(bit), .B(crc[6]), .Y(N_94_i));
    GND GND (.Y(GND_net_1));
    SLE \CRC[5]  (.D(crc[4]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[5]));
    SLE \CRC[2]  (.D(crc[1]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[2]));
    CFG2 #( .INIT(4'h6) )  \CRC_RNO[3]  (.A(N_94_i), .B(crc[2]), .Y(
        N_110_i_i));
    VCC VCC (.Y(VCC_net_1));
    SLE \CRC[4]  (.D(crc[3]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[4]));
    SLE \CRC[3]  (.D(N_110_i_i), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[3]));
    SLE \CRC[0]  (.D(N_94_i), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc[0]));
    
endmodule


module spdif_tx(
       source_right,
       source_left,
       dop_right,
       dop_left,
       reset_n_i_2,
       i2s_start,
       reset_n_i_0_RNIOUJE,
       olrck_o,
       olrck1,
       olrck2,
       use_dsd,
       spdif_tx_c,
       reset_n_i_i,
       spdif_clock_0
    );
input  [31:8] source_right;
input  [31:8] source_left;
input  [15:0] dop_right;
input  [15:0] dop_left;
output reset_n_i_2;
input  i2s_start;
input  reset_n_i_0_RNIOUJE;
output olrck_o;
input  olrck1;
input  olrck2;
input  use_dsd;
output spdif_tx_c;
input  reset_n_i_i;
input  spdif_clock_0;

    wire \bit_counter[0]_net_1 , \bit_counter_s[0] , 
        \data_out_buffer[0]_net_1 , VCC_net_1, spdif_clock_1, 
        \data_out_buffer_14[0] , GND_net_1, \data_out_buffer[1]_net_1 , 
        \data_out_buffer_14_0_iv_i[1]_net_1 , 
        \data_out_buffer[2]_net_1 , 
        \data_out_buffer_14_0_iv_i[2]_net_1 , 
        \data_out_buffer[3]_net_1 , 
        \data_out_buffer_14_0_iv_i[3]_net_1 , 
        \data_out_buffer[4]_net_1 , 
        \data_out_buffer_14_0_iv_i[4]_net_1 , 
        \data_out_buffer[5]_net_1 , 
        \data_out_buffer_14_1_iv_i[5]_net_1 , 
        \data_out_buffer[6]_net_1 , \data_out_buffer_14[6] , 
        \data_out_buffer[7]_net_1 , \data_out_buffer_14[7] , 
        \din[9]_net_1 , \din_7[9] , xsel_lr6, \din[10]_net_1 , 
        \din_7_3_i_m2_0_wmux_0_Y[10] , \din[11]_net_1 , \din_7[11] , 
        \din[12]_net_1 , \din_7_3_i_m2_0_wmux_0_Y[12] , 
        \din[13]_net_1 , \din_7[13] , \din[14]_net_1 , 
        \din_7_3_i_m2_0_wmux_0_Y[14] , \din[15]_net_1 , \din_7[15] , 
        \din[16]_net_1 , \din_7[16] , \din[17]_net_1 , \din_7[17] , 
        \din[18]_net_1 , \din_7[18] , \din[19]_net_1 , \din_7[19] , 
        \din[20]_net_1 , \din_7[20] , \din[21]_net_1 , \din_7[21] , 
        \din[22]_net_1 , \din_7[22] , \din[23]_net_1 , \din_7[23] , 
        \channel_status_shift[18]_net_1 , 
        \channel_status_shift_5[18]_net_1 , un1_frame_counter15_i, 
        \channel_status_shift[19]_net_1 , 
        \channel_status_shift_5[19]_net_1 , 
        \channel_status_shift[20]_net_1 , 
        \channel_status_shift_5[20]_net_1 , 
        \channel_status_shift[21]_net_1 , 
        \channel_status_shift_5[21]_net_1 , 
        \channel_status_shift[22]_net_1 , 
        \channel_status_shift_5[22]_net_1 , 
        \channel_status_shift[23]_net_1 , 
        \channel_status_shift_5[23]_net_1 , \din[0]_net_1 , \din_7[0] , 
        \din[1]_net_1 , \din_7[1] , \din[2]_net_1 , \din_7[2] , 
        \din[3]_net_1 , \din_7[3] , \din[4]_net_1 , \din_7[4] , 
        \din[5]_net_1 , \din_7[5] , \din[6]_net_1 , \din_7[6] , 
        \din[7]_net_1 , \din_7[7] , \din[8]_net_1 , \din_7[8] , 
        \frame_counter[6]_net_1 , un5_frame_counter_1_cry_6_S, 
        frame_counter14, \frame_counter[7]_net_1 , 
        \frame_counter_3[7]_net_1 , \frame_counter[8]_net_1 , 
        \frame_counter_3[8]_net_1 , \channel_status_shift[6]_net_1 , 
        frame_counter10_net_1, \channel_status_shift[7]_net_1 , 
        \channel_status_shift_5[7]_net_1 , 
        \channel_status_shift[8]_net_1 , 
        \channel_status_shift_5[8]_net_1 , 
        \channel_status_shift[9]_net_1 , 
        \channel_status_shift_5[9]_net_1 , 
        \channel_status_shift[10]_net_1 , 
        \channel_status_shift_5[10]_net_1 , 
        \channel_status_shift[11]_net_1 , 
        \channel_status_shift_5[11]_net_1 , 
        \channel_status_shift[12]_net_1 , 
        \channel_status_shift_5[12]_net_1 , 
        \channel_status_shift[13]_net_1 , 
        \channel_status_shift_5[13]_net_1 , 
        \channel_status_shift[14]_net_1 , 
        \channel_status_shift_5[14]_net_1 , 
        \channel_status_shift[15]_net_1 , 
        \channel_status_shift_5[15]_net_1 , 
        \channel_status_shift[16]_net_1 , 
        \channel_status_shift_5[16]_net_1 , 
        \channel_status_shift[17]_net_1 , 
        \channel_status_shift_5[17]_net_1 , \frame_counter[0]_net_1 , 
        frame_counter_96_net_1, \frame_counter[1]_net_1 , 
        un5_frame_counter_1_cry_1_S, \frame_counter[2]_net_1 , 
        un5_frame_counter_1_cry_2_S, \frame_counter[3]_net_1 , 
        un5_frame_counter_1_cry_3_S, \frame_counter[4]_net_1 , 
        un5_frame_counter_1_cry_4_S, \frame_counter[5]_net_1 , 
        un5_frame_counter_1_cry_5_S, \dop_fill[1]_net_1 , 
        dop_fill_106_net_1, \dop_fill[0]_net_1 , dop_fill_105_net_1, 
        data_biphase_0_net_1, xsel_lr, xsel_lr_0_net_1, parity_net_1, 
        parity_2_net_1, \bit_counter[1]_net_1 , \bit_counter_s[1] , 
        \bit_counter[2]_net_1 , \bit_counter_s[2] , 
        \bit_counter[3]_net_1 , \bit_counter_s[3] , 
        \bit_counter[4]_net_1 , \bit_counter_s[4] , 
        \bit_counter[5]_net_1 , \bit_counter_s[5]_net_1 , 
        bit_counter_s_413_FCO, \bit_counter_cry[1]_net_1 , 
        \bit_counter_cry[2]_net_1 , \bit_counter_cry[3]_net_1 , 
        \bit_counter_cry[4]_net_1 , un5_frame_counter_1_s_1_418_FCO, 
        un5_frame_counter_1_cry_1_net_1, 
        un5_frame_counter_1_cry_2_net_1, 
        un5_frame_counter_1_cry_3_net_1, 
        un5_frame_counter_1_cry_4_net_1, 
        un5_frame_counter_1_cry_5_net_1, 
        un5_frame_counter_1_cry_6_net_1, un5_frame_counter_1_s_8_S, 
        un5_frame_counter_1_cry_7_net_1, un5_frame_counter_1_cry_7_S, 
        \din_7_3_0_0_y0[9] , \din_7_3_0_0_co0[9] , 
        \din_7_3_0_0_y0[11] , \din_7_3_0_0_co0[11] , 
        \din_7_3_0_0_y0[2] , \din_7_3_0_0_co0[2] , \din_7_3_0_0_y0[4] , 
        \din_7_3_0_0_co0[4] , \din_7_3_0_0_y0[13] , 
        \din_7_3_0_0_co0[13] , \din_7_3_0_0_y0[15] , 
        \din_7_3_0_0_co0[15] , \din_7_3_i_m2_0_0_y0[10] , 
        \din_7_3_i_m2_0_0_co0[10] , \din_7_3_0_0_y0[8] , 
        \din_7_3_0_0_co0[8] , \din_7_3_0_0_y0[0] , 
        \din_7_3_0_0_co0[0] , \din_7_3_0_0_y0[1] , 
        \din_7_3_0_0_co0[1] , \din_7_3_0_0_y0[3] , 
        \din_7_3_0_0_co0[3] , \din_7_3_0_0_y0[7] , 
        \din_7_3_0_0_co0[7] , \din_7_3_0_0_y0[5] , 
        \din_7_3_0_0_co0[5] , \din_7_3_0_0_y0[6] , 
        \din_7_3_0_0_co0[6] , \din_7_3_i_m2_0_0_y0[12] , 
        \din_7_3_i_m2_0_0_co0[12] , \din_7_3_i_m2_0_0_y0[14] , 
        \din_7_3_i_m2_0_0_co0[14] , 
        \data_out_buffer_14_0_iv_3[0]_net_1 , 
        \data_out_buffer_14_0_iv_5[0]_net_1 , N_115_i, 
        data_out_buffer_0_sqmuxa, data_out_buffer_4_sqmuxa, 
        din_7_3_2_net_1, \din_7_3_1[16]_net_1 , din_7_3_1_net_1, 
        din_7_3_6, din_7_3_5, \din_7_3_1[23]_net_1 , 
        \din_7_3_1[22]_net_1 , \din_7_3_1[17]_net_1 , 
        \din_7_3_1[19]_net_1 , \din_7_3_1[18]_net_1 , 
        \din_7_3_1[20]_net_1 , \din_7_3_1[21]_net_1 , parity_2_6_net_1, 
        xsel_lr6_0_a2_1_net_1, N_117, \data_out_buffer_i_m[2] , 
        parity_2_17_net_1, parity_2_16_net_1, parity_2_14_net_1, 
        parity_2_13_net_1, parity_2_12_net_1, frame_counter10_5_net_1, 
        frame_counter10_4_net_1, data_out_buffer_2_sqmuxa, 
        data_out_buffer_6_sqmuxa, \data_out_buffer_14_0_iv_0[4]_net_1 , 
        parity_2_20_net_1, dop_fill_8_0_a2_3_net_1, \din_m[0] , 
        data_out_buffer_5_sqmuxa, data_out_buffer_3_sqmuxa, 
        data_out_buffer_1_sqmuxa, \din_m[19] , 
        \data_out_buffer_14_0_iv_1[2]_net_1 , 
        \data_out_buffer_14_0_iv_0[2]_net_1 , 
        \data_out_buffer_14_0_iv_1[0]_net_1 , 
        \data_out_buffer_14_0_iv_2[4]_net_1 , 
        \data_out_buffer_14_0_iv_1[6]_net_1 , parity_2_21_net_1, 
        data_out_buffer_0_sqmuxa_2_net_1, 
        \data_out_buffer_14_0_iv_4[2]_net_1 , 
        \data_out_buffer_14_0_iv_3[2]_net_1 , 
        \data_out_buffer_14_0_iv_2[2]_net_1 , 
        \data_out_buffer_14_0_iv_2[0]_net_1 , 
        \data_out_buffer_14_0_iv_4[4]_net_1 , 
        \data_out_buffer_14_0_iv_3[4]_net_1 , 
        \data_out_buffer_14_0_iv_3[6]_net_1 , 
        \data_out_buffer_14_0_iv_2[6]_net_1 ;
    
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[4]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[12]), .D(source_right[12]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[4] ), .FCO(
        \din_7_3_0_0_co0[4] ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[0]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[8]), .D(source_right[8]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[0] ), .FCO(
        \din_7_3_0_0_co0[0] ));
    SLE \channel_status_shift[18]  (.D(
        \channel_status_shift_5[18]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[18]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[8]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[7]_net_1 ), 
        .Y(\channel_status_shift_5[8]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[18]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[17]_net_1 ), 
        .Y(\channel_status_shift_5[18]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  data_out_buffer_3_sqmuxa_0_a2 (.A(
        \bit_counter[5]_net_1 ), .B(\bit_counter[4]_net_1 ), .C(
        \bit_counter[3]_net_1 ), .D(N_115_i), .Y(
        data_out_buffer_3_sqmuxa));
    SLE \channel_status_shift[16]  (.D(
        \channel_status_shift_5[16]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[16]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[23]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[22]_net_1 ), 
        .Y(\channel_status_shift_5[23]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \frame_counter_3[7]  (.A(
        frame_counter10_net_1), .B(un5_frame_counter_1_cry_7_S), .Y(
        \frame_counter_3[7]_net_1 ));
    SLE \bit_counter[3]  (.D(\bit_counter_s[3] ), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit_counter[3]_net_1 ));
    SLE \din[9]  (.D(\din_7[9] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[9]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[14]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[13]_net_1 ), 
        .Y(\channel_status_shift_5[14]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \frame_counter_3[8]  (.A(
        frame_counter10_net_1), .B(un5_frame_counter_1_s_8_S), .Y(
        \frame_counter_3[8]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  xsel_lr6_0_a2 (.A(xsel_lr6_0_a2_1_net_1)
        , .B(N_117), .C(\bit_counter[1]_net_1 ), .D(
        \bit_counter[0]_net_1 ), .Y(xsel_lr6));
    CFG4 #( .INIT(16'hFCFD) )  \din_7_3[21]  (.A(use_dsd), .B(
        din_7_3_6), .C(din_7_3_5), .D(\din_7_3_1[21]_net_1 ), .Y(
        \din_7[21] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_buffer_14_0_iv_3[0]  (.A(
        \din[23]_net_1 ), .B(\din[15]_net_1 ), .C(
        data_out_buffer_5_sqmuxa), .D(data_out_buffer_3_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_3[0]_net_1 ));
    SLE \data_out_buffer[6]  (.D(\data_out_buffer_14[6] ), .CLK(
        spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \bit_counter_s[5]  (.A(VCC_net_1), .B(
        \bit_counter[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \bit_counter_cry[4]_net_1 ), .S(\bit_counter_s[5]_net_1 ), .Y()
        , .FCO());
    SLE \channel_status_shift[10]  (.D(
        \channel_status_shift_5[10]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[10]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  frame_counter14_0_a2 (.A(
        \bit_counter[5]_net_1 ), .B(\bit_counter[4]_net_1 ), .C(
        \bit_counter[3]_net_1 ), .D(N_115_i), .Y(frame_counter14));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[0]  (.A(
        \din_7_3_0_0_y0[0] ), .B(use_dsd), .C(dop_left[0]), .D(
        dop_right[0]), .FCI(\din_7_3_0_0_co0[0] ), .S(), .Y(\din_7[0] )
        , .FCO());
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[6]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[14]), .D(source_right[14]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[6] ), .FCO(
        \din_7_3_0_0_co0[6] ));
    CFG4 #( .INIT(16'h6996) )  parity_2 (.A(parity_2_14_net_1), .B(
        parity_2_13_net_1), .C(parity_2_21_net_1), .D(
        parity_2_20_net_1), .Y(parity_2_net_1));
    SLE \din[20]  (.D(\din_7[20] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[20]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  olrck (.A(use_dsd), .B(olrck2), .C(olrck1), 
        .Y(olrck_o));
    ARI1 #( .INIT(20'h4AA00) )  \bit_counter_cry[1]  (.A(VCC_net_1), 
        .B(\bit_counter[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        bit_counter_s_413_FCO), .S(\bit_counter_s[1] ), .Y(), .FCO(
        \bit_counter_cry[1]_net_1 ));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[20]  (.A(source_left[28]), .B(
        xsel_lr), .C(source_right[28]), .Y(\din_7_3_1[20]_net_1 ));
    SLE \frame_counter[4]  (.D(un5_frame_counter_1_cry_4_S), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[4]_net_1 ));
    SLE \din[7]  (.D(\din_7[7] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[7]_net_1 ));
    SLE \bit_counter[4]  (.D(\bit_counter_s[4] ), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit_counter[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_5 (.A(
        VCC_net_1), .B(\frame_counter[5]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_cry_4_net_1), .S(
        un5_frame_counter_1_cry_5_S), .Y(), .FCO(
        un5_frame_counter_1_cry_5_net_1));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[7]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[6]_net_1 ), 
        .Y(\channel_status_shift_5[7]_net_1 ));
    CFG3 #( .INIT(8'hBA) )  \data_out_buffer_14_0_iv_3[2]  (.A(
        \data_out_buffer_14_0_iv_1[2]_net_1 ), .B(\din[22]_net_1 ), .C(
        data_out_buffer_5_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_3[2]_net_1 ));
    CFG4 #( .INIT(16'hFFF2) )  \data_out_buffer_14_0_iv_2[6]  (.A(
        \data_out_buffer[5]_net_1 ), .B(N_115_i), .C(\din_m[0] ), .D(
        \data_out_buffer_14_0_iv_1[6]_net_1 ), .Y(
        \data_out_buffer_14_0_iv_2[6]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  data_out_buffer_1_sqmuxa_0_a2 (.A(
        \bit_counter[5]_net_1 ), .B(\bit_counter[4]_net_1 ), .C(
        \bit_counter[3]_net_1 ), .D(N_115_i), .Y(
        data_out_buffer_1_sqmuxa));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[9]  (.A(
        \din_7_3_0_0_y0[9] ), .B(use_dsd), .C(dop_left[9]), .D(
        dop_right[9]), .FCI(\din_7_3_0_0_co0[9] ), .S(), .Y(\din_7[9] )
        , .FCO());
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[2]  (.A(
        \din_7_3_0_0_y0[2] ), .B(use_dsd), .C(dop_left[2]), .D(
        dop_right[2]), .FCI(\din_7_3_0_0_co0[2] ), .S(), .Y(\din_7[2] )
        , .FCO());
    CFG4 #( .INIT(16'h0023) )  \data_out_buffer_14_0_iv_i[3]  (.A(
        \frame_counter[0]_net_1 ), .B(\data_out_buffer_i_m[2] ), .C(
        frame_counter14), .D(data_out_buffer_0_sqmuxa_2_net_1), .Y(
        \data_out_buffer_14_0_iv_i[3]_net_1 ));
    CFG3 #( .INIT(8'hBA) )  \data_out_buffer_14_0_iv_2[2]  (.A(
        \data_out_buffer_14_0_iv_0[2]_net_1 ), .B(\din[2]_net_1 ), .C(
        data_out_buffer_0_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_2[2]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  parity_2_14 (.A(\din[6]_net_1 ), .B(
        \din[5]_net_1 ), .C(\din[4]_net_1 ), .D(\din[3]_net_1 ), .Y(
        parity_2_14_net_1));
    SLE \frame_counter[1]  (.D(un5_frame_counter_1_cry_1_S), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_s_1_418 (.A(
        VCC_net_1), .B(\frame_counter[0]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        un5_frame_counter_1_s_1_418_FCO));
    CLKINT spdif_clock_1_RNO (.A(spdif_clock_0), .Y(spdif_clock_1));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_2 (.A(
        VCC_net_1), .B(\frame_counter[2]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_cry_1_net_1), .S(
        un5_frame_counter_1_cry_2_S), .Y(), .FCO(
        un5_frame_counter_1_cry_2_net_1));
    CFG4 #( .INIT(16'hFEEE) )  \data_out_buffer_14_0_iv[0]  (.A(
        \data_out_buffer_14_0_iv_2[0]_net_1 ), .B(
        \data_out_buffer_14_0_iv_5[0]_net_1 ), .C(\din[7]_net_1 ), .D(
        data_out_buffer_1_sqmuxa), .Y(\data_out_buffer_14[0] ));
    GND GND (.Y(GND_net_1));
    SLE \din[5]  (.D(\din_7[5] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[5]_net_1 ));
    CFG3 #( .INIT(8'h20) )  din_7_3_13 (.A(\dop_fill[1]_net_1 ), .B(
        xsel_lr), .C(use_dsd), .Y(din_7_3_5));
    SLE \channel_status_shift[19]  (.D(
        \channel_status_shift_5[19]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[19]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  data_out_buffer_4_sqmuxa_0_a2 (.A(
        \bit_counter[4]_net_1 ), .B(\bit_counter[3]_net_1 ), .C(
        N_115_i), .D(\bit_counter[5]_net_1 ), .Y(
        data_out_buffer_4_sqmuxa));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[4]  (.A(
        \din_7_3_0_0_y0[4] ), .B(use_dsd), .C(dop_left[4]), .D(
        dop_right[4]), .FCI(\din_7_3_0_0_co0[4] ), .S(), .Y(\din_7[4] )
        , .FCO());
    SLE \data_out_buffer[4]  (.D(\data_out_buffer_14_0_iv_i[4]_net_1 ), 
        .CLK(spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[4]_net_1 ));
    SLE \channel_status_shift[6]  (.D(frame_counter10_net_1), .CLK(
        spdif_clock_1), .EN(un1_frame_counter15_i), .ALn(reset_n_i_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\channel_status_shift[6]_net_1 ));
    SLE \frame_counter[2]  (.D(un5_frame_counter_1_cry_2_S), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[16]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[15]_net_1 ), 
        .Y(\channel_status_shift_5[16]_net_1 ));
    SLE \data_out_buffer[3]  (.D(\data_out_buffer_14_0_iv_i[3]_net_1 ), 
        .CLK(spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[3]_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  \data_out_buffer_14_0_iv_3[4]  (.A(
        \data_out_buffer_14_0_iv_0[4]_net_1 ), .B(
        \data_out_buffer_14_0_iv_2[4]_net_1 ), .C(\din[17]_net_1 ), .D(
        data_out_buffer_4_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_3[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \data_out_buffer_14_0_iv_2_RNO[6]  (.A(
        data_out_buffer_0_sqmuxa), .B(\din[0]_net_1 ), .Y(\din_m[0] ));
    CFG4 #( .INIT(16'hFCFD) )  \din_7_3[23]  (.A(use_dsd), .B(
        din_7_3_6), .C(din_7_3_5), .D(\din_7_3_1[23]_net_1 ), .Y(
        \din_7[23] ));
    SLE \din[15]  (.D(\din_7[15] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[15]_net_1 ));
    SLE \channel_status_shift[7]  (.D(
        \channel_status_shift_5[7]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[7]_net_1 ));
    CFG2 #( .INIT(4'h6) )  xsel_lr_0 (.A(xsel_lr6), .B(xsel_lr), .Y(
        xsel_lr_0_net_1));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[17]  (.A(source_left[25]), .B(
        xsel_lr), .C(source_right[25]), .Y(\din_7_3_1[17]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  frame_counter10_5 (.A(
        \frame_counter[8]_net_1 ), .B(\frame_counter[6]_net_1 ), .C(
        \frame_counter[5]_net_1 ), .D(\frame_counter[4]_net_1 ), .Y(
        frame_counter10_5_net_1));
    CFG3 #( .INIT(8'h20) )  din_7_3_1 (.A(\dop_fill[0]_net_1 ), .B(
        xsel_lr), .C(use_dsd), .Y(din_7_3_1_net_1));
    SLE \frame_counter[6]  (.D(un5_frame_counter_1_cry_6_S), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[6]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[5]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[13]), .D(source_right[13]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[5] ), .FCO(
        \din_7_3_0_0_co0[5] ));
    CFG4 #( .INIT(16'h0EEE) )  \data_out_buffer_14_0_iv_i[1]  (.A(
        N_115_i), .B(\data_out_buffer[0]_net_1 ), .C(frame_counter14), 
        .D(frame_counter10_net_1), .Y(
        \data_out_buffer_14_0_iv_i[1]_net_1 ));
    SLE \data_out_buffer[0]  (.D(\data_out_buffer_14[0] ), .CLK(
        spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[17]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[16]_net_1 ), 
        .Y(\channel_status_shift_5[17]_net_1 ));
    SLE \channel_status_shift[21]  (.D(
        \channel_status_shift_5[21]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[21]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_i_m2_0_0_wmux[10]  (.A(
        xsel_lr), .B(use_dsd), .C(source_left[18]), .D(
        source_right[18]), .FCI(VCC_net_1), .S(), .Y(
        \din_7_3_i_m2_0_0_y0[10] ), .FCO(\din_7_3_i_m2_0_0_co0[10] ));
    SLE \channel_status_shift[22]  (.D(
        \channel_status_shift_5[22]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[22]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  parity_2_20 (.A(\din[7]_net_1 ), .B(
        \din[8]_net_1 ), .C(parity_2_16_net_1), .D(parity_2_6_net_1), 
        .Y(parity_2_20_net_1));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[8]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[16]), .D(source_right[16]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[8] ), .FCO(
        \din_7_3_0_0_co0[8] ));
    CFG4 #( .INIT(16'h0001) )  \data_out_buffer_14_0_iv_i[2]  (.A(
        \data_out_buffer_14_0_iv_2[2]_net_1 ), .B(
        \data_out_buffer_14_0_iv_3[2]_net_1 ), .C(
        \data_out_buffer_14_0_iv_4[2]_net_1 ), .D(
        data_out_buffer_0_sqmuxa_2_net_1), .Y(
        \data_out_buffer_14_0_iv_i[2]_net_1 ));
    SLE \din[16]  (.D(\din_7[16] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[16]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \data_out_buffer_14_0_iv_2_RNO[0]  (.A(
        data_out_buffer_4_sqmuxa), .B(\din[19]_net_1 ), .Y(\din_m[19] )
        );
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_6 (.A(
        VCC_net_1), .B(\frame_counter[6]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_cry_5_net_1), .S(
        un5_frame_counter_1_cry_6_S), .Y(), .FCO(
        un5_frame_counter_1_cry_6_net_1));
    SLE \data_out_buffer[2]  (.D(\data_out_buffer_14_0_iv_i[2]_net_1 ), 
        .CLK(spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[2]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \data_out_buffer_14_0_iv_1[2]  (.A(
        \din[18]_net_1 ), .B(\din[10]_net_1 ), .C(
        data_out_buffer_4_sqmuxa), .D(data_out_buffer_2_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_1[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[22]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[21]_net_1 ), 
        .Y(\channel_status_shift_5[22]_net_1 ));
    SLE \din[3]  (.D(\din_7[3] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[3]_net_1 ));
    SLE data_biphase (.D(data_biphase_0_net_1), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(spdif_tx_c));
    SLE \bit_counter[2]  (.D(\bit_counter_s[2] ), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit_counter[2]_net_1 ));
    SLE \frame_counter[0]  (.D(frame_counter_96_net_1), .CLK(
        spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[11]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[10]_net_1 ), 
        .Y(\channel_status_shift_5[11]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_4 (.A(
        VCC_net_1), .B(\frame_counter[4]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_cry_3_net_1), .S(
        un5_frame_counter_1_cry_4_S), .Y(), .FCO(
        un5_frame_counter_1_cry_4_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_1 (.A(
        VCC_net_1), .B(\frame_counter[1]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_s_1_418_FCO), .S(
        un5_frame_counter_1_cry_1_S), .Y(), .FCO(
        un5_frame_counter_1_cry_1_net_1));
    SLE \channel_status_shift[23]  (.D(
        \channel_status_shift_5[23]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[23]_net_1 ));
    SLE \channel_status_shift[8]  (.D(
        \channel_status_shift_5[8]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[8]_net_1 ));
    CFG3 #( .INIT(8'h96) )  parity_2_12 (.A(\din[23]_net_1 ), .B(
        \din[22]_net_1 ), .C(\din[21]_net_1 ), .Y(parity_2_12_net_1));
    SLE \data_out_buffer[7]  (.D(\data_out_buffer_14[7] ), .CLK(
        spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[7]_net_1 ));
    CFG4 #( .INIT(16'hF870) )  dop_fill_105 (.A(N_117), .B(
        dop_fill_8_0_a2_3_net_1), .C(\dop_fill[0]_net_1 ), .D(
        \dop_fill[1]_net_1 ), .Y(dop_fill_105_net_1));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_i_m2_0_wmux_0[14]  (.A(
        \din_7_3_i_m2_0_0_y0[14] ), .B(use_dsd), .C(dop_left[14]), .D(
        dop_right[14]), .FCI(\din_7_3_i_m2_0_0_co0[14] ), .S(), .Y(
        \din_7_3_i_m2_0_wmux_0_Y[14] ), .FCO());
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[15]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[14]_net_1 ), 
        .Y(\channel_status_shift_5[15]_net_1 ));
    SLE \din[11]  (.D(\din_7[11] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[11]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[6]  (.A(
        \din_7_3_0_0_y0[6] ), .B(use_dsd), .C(dop_left[6]), .D(
        dop_right[6]), .FCI(\din_7_3_0_0_co0[6] ), .S(), .Y(\din_7[6] )
        , .FCO());
    CFG3 #( .INIT(8'h08) )  data_out_buffer_0_sqmuxa_2 (.A(
        frame_counter14), .B(\frame_counter[0]_net_1 ), .C(
        frame_counter10_net_1), .Y(data_out_buffer_0_sqmuxa_2_net_1));
    SLE \frame_counter[3]  (.D(un5_frame_counter_1_cry_3_S), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[3]_net_1 ));
    SLE \din[8]  (.D(\din_7[8] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[8]_net_1 ));
    SLE \din[18]  (.D(\din_7[18] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[18]_net_1 ));
    SLE \data_out_buffer[5]  (.D(\data_out_buffer_14_1_iv_i[5]_net_1 ), 
        .CLK(spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[5]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[1]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[9]), .D(source_right[9]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[1] ), .FCO(
        \din_7_3_0_0_co0[1] ));
    CFG3 #( .INIT(8'h80) )  data_out_buffer65_i_a2 (.A(
        \bit_counter[2]_net_1 ), .B(\bit_counter[1]_net_1 ), .C(
        \bit_counter[0]_net_1 ), .Y(N_115_i));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_i_m2_0_0_wmux[12]  (.A(
        xsel_lr), .B(use_dsd), .C(source_left[20]), .D(
        source_right[20]), .FCI(VCC_net_1), .S(), .Y(
        \din_7_3_i_m2_0_0_y0[12] ), .FCO(\din_7_3_i_m2_0_0_co0[12] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_buffer_14_0_iv_1[6]  (.A(
        \din[16]_net_1 ), .B(\din[8]_net_1 ), .C(
        data_out_buffer_4_sqmuxa), .D(data_out_buffer_2_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_1[6]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[3]  (.A(
        \din_7_3_0_0_y0[3] ), .B(use_dsd), .C(dop_left[3]), .D(
        dop_right[3]), .FCI(\din_7_3_0_0_co0[3] ), .S(), .Y(\din_7[3] )
        , .FCO());
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[10]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[9]_net_1 ), 
        .Y(\channel_status_shift_5[10]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  data_out_buffer_2_sqmuxa_0_a2 (.A(
        \bit_counter[5]_net_1 ), .B(\bit_counter[4]_net_1 ), .C(
        \bit_counter[3]_net_1 ), .D(N_115_i), .Y(
        data_out_buffer_2_sqmuxa));
    CFG4 #( .INIT(16'hECA0) )  \data_out_buffer_14_0_iv_3[6]  (.A(
        \din[20]_net_1 ), .B(\din[12]_net_1 ), .C(
        data_out_buffer_5_sqmuxa), .D(data_out_buffer_3_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_3[6]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  frame_counter10 (.A(
        \frame_counter[7]_net_1 ), .B(\frame_counter[1]_net_1 ), .C(
        frame_counter10_5_net_1), .D(frame_counter10_4_net_1), .Y(
        frame_counter10_net_1));
    SLE \din[14]  (.D(\din_7_3_i_m2_0_wmux_0_Y[14] ), .CLK(
        spdif_clock_1), .EN(xsel_lr6), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\din[14]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[7]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[15]), .D(source_right[15]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[7] ), .FCO(
        \din_7_3_0_0_co0[7] ));
    CFG4 #( .INIT(16'h6996) )  parity_2_17 (.A(\din[18]_net_1 ), .B(
        \din[17]_net_1 ), .C(\din[16]_net_1 ), .D(\din[15]_net_1 ), .Y(
        parity_2_17_net_1));
    CFG2 #( .INIT(4'h1) )  xsel_lr6_0_a2_0 (.A(\bit_counter[3]_net_1 ), 
        .B(\bit_counter[4]_net_1 ), .Y(N_117));
    CFG3 #( .INIT(8'h80) )  din_7_3_2 (.A(\dop_fill[0]_net_1 ), .B(
        xsel_lr), .C(use_dsd), .Y(din_7_3_2_net_1));
    CFG4 #( .INIT(16'h05CD) )  \data_out_buffer_14_0_iv_0[2]  (.A(
        N_115_i), .B(data_out_buffer_6_sqmuxa), .C(
        \data_out_buffer[1]_net_1 ), .D(
        \channel_status_shift[23]_net_1 ), .Y(
        \data_out_buffer_14_0_iv_0[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[13]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[12]_net_1 ), 
        .Y(\channel_status_shift_5[13]_net_1 ));
    SLE \din[21]  (.D(\din_7[21] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[21]_net_1 ));
    SLE \dop_fill[0]  (.D(dop_fill_105_net_1), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dop_fill[0]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[15]  (.A(xsel_lr), 
        .B(use_dsd), .C(source_left[23]), .D(source_right[23]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[15] ), .FCO(
        \din_7_3_0_0_co0[15] ));
    SLE \frame_counter[5]  (.D(un5_frame_counter_1_cry_5_S), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[5]_net_1 ));
    SLE \channel_status_shift[20]  (.D(
        \channel_status_shift_5[20]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[20]_net_1 ));
    CFG3 #( .INIT(8'h80) )  frame_counter10_4 (.A(
        \frame_counter[3]_net_1 ), .B(\frame_counter[2]_net_1 ), .C(
        \frame_counter[0]_net_1 ), .Y(frame_counter10_4_net_1));
    SLE \frame_counter[7]  (.D(\frame_counter_3[7]_net_1 ), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[7]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  data_out_buffer_6_sqmuxa_0_a2 (.A(
        \bit_counter[5]_net_1 ), .B(\bit_counter[4]_net_1 ), .C(
        \bit_counter[3]_net_1 ), .D(N_115_i), .Y(
        data_out_buffer_6_sqmuxa));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[2]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[10]), .D(source_right[10]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[2] ), .FCO(
        \din_7_3_0_0_co0[2] ));
    CFG3 #( .INIT(8'h32) )  \data_out_buffer_14_1_iv_i[5]  (.A(N_115_i)
        , .B(frame_counter14), .C(\data_out_buffer[4]_net_1 ), .Y(
        \data_out_buffer_14_1_iv_i[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \bit_counter_cry[2]  (.A(VCC_net_1), 
        .B(\bit_counter[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \bit_counter_cry[1]_net_1 ), .S(\bit_counter_s[2] ), .Y(), 
        .FCO(\bit_counter_cry[2]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  parity_2_21 (.A(\din[19]_net_1 ), .B(
        \din[20]_net_1 ), .C(parity_2_17_net_1), .D(parity_2_12_net_1), 
        .Y(parity_2_21_net_1));
    SLE parity (.D(parity_2_net_1), .CLK(spdif_clock_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(parity_net_1));
    SLE \din[2]  (.D(\din_7[2] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \bit_counter_RNO[0]  (.A(
        \bit_counter[0]_net_1 ), .Y(\bit_counter_s[0] ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[13]  (.A(xsel_lr), 
        .B(use_dsd), .C(source_left[21]), .D(source_right[21]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[13] ), .FCO(
        \din_7_3_0_0_co0[13] ));
    ARI1 #( .INIT(20'h4AA00) )  \bit_counter_cry[3]  (.A(VCC_net_1), 
        .B(\bit_counter[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \bit_counter_cry[2]_net_1 ), .S(\bit_counter_s[3] ), .Y(), 
        .FCO(\bit_counter_cry[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[9]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[8]_net_1 ), 
        .Y(\channel_status_shift_5[9]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[13]  (.A(
        \din_7_3_0_0_y0[13] ), .B(use_dsd), .C(dop_left[13]), .D(
        dop_right[13]), .FCI(\din_7_3_0_0_co0[13] ), .S(), .Y(
        \din_7[13] ), .FCO());
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[8]  (.A(
        \din_7_3_0_0_y0[8] ), .B(use_dsd), .C(dop_left[8]), .D(
        dop_right[8]), .FCI(\din_7_3_0_0_co0[8] ), .S(), .Y(\din_7[8] )
        , .FCO());
    CFG3 #( .INIT(8'hCD) )  \data_out_buffer_14_0_iv_0[4]  (.A(N_115_i)
        , .B(data_out_buffer_6_sqmuxa), .C(\data_out_buffer[3]_net_1 ), 
        .Y(\data_out_buffer_14_0_iv_0[4]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_i_m2_0_wmux_0[10]  (.A(
        \din_7_3_i_m2_0_0_y0[10] ), .B(use_dsd), .C(dop_left[10]), .D(
        dop_right[10]), .FCI(\din_7_3_i_m2_0_0_co0[10] ), .S(), .Y(
        \din_7_3_i_m2_0_wmux_0_Y[10] ), .FCO());
    CFG2 #( .INIT(4'hE) )  \data_out_buffer_RNO[7]  (.A(N_115_i), .B(
        \data_out_buffer[6]_net_1 ), .Y(\data_out_buffer_14[7] ));
    CFG2 #( .INIT(4'h6) )  data_biphase_0 (.A(spdif_tx_c), .B(
        \data_out_buffer[7]_net_1 ), .Y(data_biphase_0_net_1));
    CFG3 #( .INIT(8'h80) )  din_7_3_10 (.A(\dop_fill[1]_net_1 ), .B(
        xsel_lr), .C(use_dsd), .Y(din_7_3_6));
    SLE \din[19]  (.D(\din_7[19] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  bit_counter_s_413 (.A(VCC_net_1), .B(
        \bit_counter[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(bit_counter_s_413_FCO));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[11]  (.A(
        \din_7_3_0_0_y0[11] ), .B(use_dsd), .C(dop_left[11]), .D(
        dop_right[11]), .FCI(\din_7_3_0_0_co0[11] ), .S(), .Y(
        \din_7[11] ), .FCO());
    CFG2 #( .INIT(4'h4) )  reset_n_i (.A(reset_n_i_0_RNIOUJE), .B(
        i2s_start), .Y(reset_n_i_2));
    CFG4 #( .INIT(16'h0020) )  dop_fill_8_0_a2_3 (.A(
        \bit_counter[0]_net_1 ), .B(\bit_counter[1]_net_1 ), .C(
        xsel_lr6_0_a2_1_net_1), .D(xsel_lr), .Y(
        dop_fill_8_0_a2_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_s_8 (.A(VCC_net_1), 
        .B(\frame_counter[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un5_frame_counter_1_cry_7_net_1), .S(
        un5_frame_counter_1_s_8_S), .Y(), .FCO());
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[22]  (.A(source_left[30]), .B(
        xsel_lr), .C(source_right[30]), .Y(\din_7_3_1[22]_net_1 ));
    CFG4 #( .INIT(16'hFFAB) )  \din_7_3[18]  (.A(din_7_3_2_net_1), .B(
        use_dsd), .C(\din_7_3_1[18]_net_1 ), .D(din_7_3_1_net_1), .Y(
        \din_7[18] ));
    SLE \frame_counter[8]  (.D(\frame_counter_3[8]_net_1 ), .CLK(
        spdif_clock_1), .EN(frame_counter14), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\frame_counter[8]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[3]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[11]), .D(source_right[11]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[3] ), .FCO(
        \din_7_3_0_0_co0[3] ));
    CFG4 #( .INIT(16'hFCFD) )  \din_7_3[20]  (.A(use_dsd), .B(
        din_7_3_6), .C(din_7_3_5), .D(\din_7_3_1[20]_net_1 ), .Y(
        \din_7[20] ));
    SLE xsel_lr_1 (.D(xsel_lr_0_net_1), .CLK(spdif_clock_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(xsel_lr));
    CFG2 #( .INIT(4'h6) )  parity_2_6 (.A(\din[9]_net_1 ), .B(
        \din[10]_net_1 ), .Y(parity_2_6_net_1));
    SLE \din[13]  (.D(\din_7[13] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[13]_net_1 ));
    SLE \din[17]  (.D(\din_7[17] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[17]_net_1 ));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[19]  (.A(source_left[27]), .B(
        xsel_lr), .C(source_right[27]), .Y(\din_7_3_1[19]_net_1 ));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[23]  (.A(source_left[31]), .B(
        xsel_lr), .C(source_right[31]), .Y(\din_7_3_1[23]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \data_out_buffer_14_0_iv_4[4]  (.A(
        \din[21]_net_1 ), .B(\din[13]_net_1 ), .C(
        data_out_buffer_5_sqmuxa), .D(data_out_buffer_3_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_4[4]_net_1 ));
    SLE \channel_status_shift[9]  (.D(
        \channel_status_shift_5[9]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[9]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[1]  (.A(
        \din_7_3_0_0_y0[1] ), .B(use_dsd), .C(dop_left[1]), .D(
        dop_right[1]), .FCI(\din_7_3_0_0_co0[1] ), .S(), .Y(\din_7[1] )
        , .FCO());
    SLE \din[0]  (.D(\din_7[0] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  frame_counter_96 (.A(frame_counter14), .B(
        \frame_counter[0]_net_1 ), .Y(frame_counter_96_net_1));
    SLE \din[4]  (.D(\din_7[4] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[4]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  data_out_buffer_0_sqmuxa_0_a2 (.A(
        \bit_counter[4]_net_1 ), .B(\bit_counter[3]_net_1 ), .C(
        N_115_i), .D(\bit_counter[5]_net_1 ), .Y(
        data_out_buffer_0_sqmuxa));
    CFG4 #( .INIT(16'hFFAB) )  \din_7_3[16]  (.A(din_7_3_2_net_1), .B(
        use_dsd), .C(\din_7_3_1[16]_net_1 ), .D(din_7_3_1_net_1), .Y(
        \din_7[16] ));
    CFG4 #( .INIT(16'hFCFD) )  \din_7_3[22]  (.A(use_dsd), .B(
        din_7_3_6), .C(din_7_3_5), .D(\din_7_3_1[22]_net_1 ), .Y(
        \din_7[22] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_buffer_14_0_iv_1[0]  (.A(
        \din[3]_net_1 ), .B(\din[11]_net_1 ), .C(
        data_out_buffer_2_sqmuxa), .D(data_out_buffer_0_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_1[0]_net_1 ));
    SLE \din[12]  (.D(\din_7_3_i_m2_0_wmux_0_Y[12] ), .CLK(
        spdif_clock_1), .EN(xsel_lr6), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\din[12]_net_1 ));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[21]  (.A(source_left[29]), .B(
        xsel_lr), .C(source_right[29]), .Y(\din_7_3_1[21]_net_1 ));
    SLE \bit_counter[5]  (.D(\bit_counter_s[5]_net_1 ), .CLK(
        spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\bit_counter[5]_net_1 ));
    SLE \din[1]  (.D(\din_7[1] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[1]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  \data_out_buffer_14_0_iv_2[4]  (.A(
        \din[1]_net_1 ), .B(\din[9]_net_1 ), .C(
        data_out_buffer_2_sqmuxa), .D(data_out_buffer_0_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_2[4]_net_1 ));
    SLE \din[23]  (.D(\din_7[23] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[23]_net_1 ));
    CFG4 #( .INIT(16'hF4F0) )  \data_out_buffer_14_0_iv_5[0]  (.A(
        frame_counter10_net_1), .B(\frame_counter[0]_net_1 ), .C(
        \data_out_buffer_14_0_iv_3[0]_net_1 ), .D(frame_counter14), .Y(
        \data_out_buffer_14_0_iv_5[0]_net_1 ));
    SLE \channel_status_shift[11]  (.D(
        \channel_status_shift_5[11]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[11]_net_1 ));
    SLE \channel_status_shift[12]  (.D(
        \channel_status_shift_5[12]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[12]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_i_m2_0_wmux_0[12]  (.A(
        \din_7_3_i_m2_0_0_y0[12] ), .B(use_dsd), .C(dop_left[12]), .D(
        dop_right[12]), .FCI(\din_7_3_i_m2_0_0_co0[12] ), .S(), .Y(
        \din_7_3_i_m2_0_wmux_0_Y[12] ), .FCO());
    CFG4 #( .INIT(16'h2000) )  data_out_buffer_5_sqmuxa_0_a2 (.A(
        \bit_counter[5]_net_1 ), .B(\bit_counter[4]_net_1 ), .C(
        \bit_counter[3]_net_1 ), .D(N_115_i), .Y(
        data_out_buffer_5_sqmuxa));
    CFG4 #( .INIT(16'h1011) )  \data_out_buffer_14_0_iv_i[4]  (.A(
        \data_out_buffer_14_0_iv_4[4]_net_1 ), .B(
        \data_out_buffer_14_0_iv_3[4]_net_1 ), .C(\din[5]_net_1 ), .D(
        data_out_buffer_1_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_i[4]_net_1 ));
    CFG4 #( .INIT(16'hFEEE) )  \data_out_buffer_14_0_iv[6]  (.A(
        \data_out_buffer_14_0_iv_3[6]_net_1 ), .B(
        \data_out_buffer_14_0_iv_2[6]_net_1 ), .C(\din[4]_net_1 ), .D(
        data_out_buffer_1_sqmuxa), .Y(\data_out_buffer_14[6] ));
    SLE \bit_counter[0]  (.D(\bit_counter_s[0] ), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit_counter[0]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[7]  (.A(
        \din_7_3_0_0_y0[7] ), .B(use_dsd), .C(dop_left[7]), .D(
        dop_right[7]), .FCI(\din_7_3_0_0_co0[7] ), .S(), .Y(\din_7[7] )
        , .FCO());
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[5]  (.A(
        \din_7_3_0_0_y0[5] ), .B(use_dsd), .C(dop_left[5]), .D(
        dop_right[5]), .FCI(\din_7_3_0_0_co0[5] ), .S(), .Y(\din_7[5] )
        , .FCO());
    CFG4 #( .INIT(16'hFCFD) )  \din_7_3[17]  (.A(use_dsd), .B(
        din_7_3_6), .C(din_7_3_5), .D(\din_7_3_1[17]_net_1 ), .Y(
        \din_7[17] ));
    SLE \din[22]  (.D(\din_7[22] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[22]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \data_out_buffer_14_0_iv_4[2]  (.A(
        \din[14]_net_1 ), .B(\din[6]_net_1 ), .C(
        data_out_buffer_3_sqmuxa), .D(data_out_buffer_1_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_4[2]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \channel_status_shift_5[21]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[20]_net_1 ), 
        .Y(\channel_status_shift_5[21]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  parity_2_13 (.A(\din[2]_net_1 ), .B(
        \din[1]_net_1 ), .C(\din[0]_net_1 ), .D(
        \channel_status_shift[23]_net_1 ), .Y(parity_2_13_net_1));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[18]  (.A(source_left[26]), .B(
        xsel_lr), .C(source_right[26]), .Y(\din_7_3_1[18]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[9]  (.A(xsel_lr), .B(
        use_dsd), .C(source_left[17]), .D(source_right[17]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[9] ), .FCO(
        \din_7_3_0_0_co0[9] ));
    SLE \din[6]  (.D(\din_7[6] ), .CLK(spdif_clock_1), .EN(xsel_lr6), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\din[6]_net_1 ));
    SLE \channel_status_shift[13]  (.D(
        \channel_status_shift_5[13]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[13]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_3 (.A(
        VCC_net_1), .B(\frame_counter[3]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_cry_2_net_1), .S(
        un5_frame_counter_1_cry_3_S), .Y(), .FCO(
        un5_frame_counter_1_cry_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un5_frame_counter_1_cry_7 (.A(
        VCC_net_1), .B(\frame_counter[7]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un5_frame_counter_1_cry_6_net_1), .S(
        un5_frame_counter_1_cry_7_S), .Y(), .FCO(
        un5_frame_counter_1_cry_7_net_1));
    CFG4 #( .INIT(16'h6996) )  parity_2_16 (.A(\din[14]_net_1 ), .B(
        \din[13]_net_1 ), .C(\din[12]_net_1 ), .D(\din[11]_net_1 ), .Y(
        parity_2_16_net_1));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_i_m2_0_0_wmux[14]  (.A(
        xsel_lr), .B(use_dsd), .C(source_left[22]), .D(
        source_right[22]), .FCI(VCC_net_1), .S(), .Y(
        \din_7_3_i_m2_0_0_y0[14] ), .FCO(\din_7_3_i_m2_0_0_co0[14] ));
    CFG4 #( .INIT(16'hFEEE) )  \data_out_buffer_14_0_iv_2[0]  (.A(
        \din_m[19] ), .B(\data_out_buffer_14_0_iv_1[0]_net_1 ), .C(
        parity_net_1), .D(data_out_buffer_6_sqmuxa), .Y(
        \data_out_buffer_14_0_iv_2[0]_net_1 ));
    SLE \bit_counter[1]  (.D(\bit_counter_s[1] ), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit_counter[1]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \din_7_3_0_0_wmux[11]  (.A(xsel_lr), 
        .B(use_dsd), .C(source_left[19]), .D(source_right[19]), .FCI(
        VCC_net_1), .S(), .Y(\din_7_3_0_0_y0[11] ), .FCO(
        \din_7_3_0_0_co0[11] ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[12]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[11]_net_1 ), 
        .Y(\channel_status_shift_5[12]_net_1 ));
    SLE \channel_status_shift[14]  (.D(
        \channel_status_shift_5[14]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[14]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \din_7_3_0_wmux_0[15]  (.A(
        \din_7_3_0_0_y0[15] ), .B(use_dsd), .C(dop_left[15]), .D(
        dop_right[15]), .FCI(\din_7_3_0_0_co0[15] ), .S(), .Y(
        \din_7[15] ), .FCO());
    CFG2 #( .INIT(4'h1) )  xsel_lr6_0_a2_1 (.A(\bit_counter[5]_net_1 ), 
        .B(\bit_counter[2]_net_1 ), .Y(xsel_lr6_0_a2_1_net_1));
    SLE \dop_fill[1]  (.D(dop_fill_106_net_1), .CLK(spdif_clock_1), 
        .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dop_fill[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \bit_counter_cry[4]  (.A(VCC_net_1), 
        .B(\bit_counter[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \bit_counter_cry[3]_net_1 ), .S(\bit_counter_s[4] ), .Y(), 
        .FCO(\bit_counter_cry[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \frame_counter_RNIC7RL[0]  (.A(
        frame_counter14), .B(\frame_counter[0]_net_1 ), .Y(
        un1_frame_counter15_i));
    CFG3 #( .INIT(8'h1D) )  \din_7_3_1[16]  (.A(source_left[24]), .B(
        xsel_lr), .C(source_right[24]), .Y(\din_7_3_1[16]_net_1 ));
    SLE \data_out_buffer[1]  (.D(\data_out_buffer_14_0_iv_i[1]_net_1 ), 
        .CLK(spdif_clock_1), .EN(VCC_net_1), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\data_out_buffer[1]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \data_out_buffer_14_0_iv_i_RNO[3]  (.A(
        N_115_i), .B(\data_out_buffer[2]_net_1 ), .Y(
        \data_out_buffer_i_m[2] ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[20]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[19]_net_1 ), 
        .Y(\channel_status_shift_5[20]_net_1 ));
    SLE \channel_status_shift[15]  (.D(
        \channel_status_shift_5[15]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[15]_net_1 ));
    CFG4 #( .INIT(16'hFCFD) )  \din_7_3[19]  (.A(use_dsd), .B(
        din_7_3_6), .C(din_7_3_5), .D(\din_7_3_1[19]_net_1 ), .Y(
        \din_7[19] ));
    CFG2 #( .INIT(4'h4) )  \channel_status_shift_5[19]  (.A(
        frame_counter10_net_1), .B(\channel_status_shift[18]_net_1 ), 
        .Y(\channel_status_shift_5[19]_net_1 ));
    SLE \din[10]  (.D(\din_7_3_i_m2_0_wmux_0_Y[10] ), .CLK(
        spdif_clock_1), .EN(xsel_lr6), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\din[10]_net_1 ));
    SLE \channel_status_shift[17]  (.D(
        \channel_status_shift_5[17]_net_1 ), .CLK(spdif_clock_1), .EN(
        un1_frame_counter15_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \channel_status_shift[17]_net_1 ));
    CFG3 #( .INIT(8'h78) )  dop_fill_106 (.A(N_117), .B(
        dop_fill_8_0_a2_3_net_1), .C(\dop_fill[1]_net_1 ), .Y(
        dop_fill_106_net_1));
    
endmodule


module sync_logic_1s_1(
       sound_card_ctrl_0,
       sdctrl_use_dsd,
       sdclk_n_1,
       mclk_1,
       N_4047_i
    );
input  sound_card_ctrl_0;
output sdctrl_use_dsd;
input  sdclk_n_1;
input  mclk_1;
input  N_4047_i;

    wire \update_ack_dly[1]_net_1 , \update_ack_dly_i[1] , 
        \update_strobe_dly[1]_net_1 , VCC_net_1, 
        \update_strobe_dly[0]_net_1 , GND_net_1, 
        \update_strobe_dly[2]_net_1 , \update_strobe_dly[3]_net_1 , 
        update_strobe_net_1, update_ack_net_1, \data_buf[0]_net_1 , 
        un1_update_strobe_dly_0, data_buf6_i_net_1, 
        \update_ack_dly[0]_net_1 ;
    
    SLE update_strobe (.D(\update_ack_dly_i[1] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(update_strobe_net_1));
    GND GND (.Y(GND_net_1));
    SLE \data_buf_sync[0]  (.D(\data_buf[0]_net_1 ), .CLK(mclk_1), .EN(
        un1_update_strobe_dly_0), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdctrl_use_dsd));
    CFG2 #( .INIT(4'h9) )  data_buf6_i (.A(update_strobe_net_1), .B(
        \update_ack_dly[1]_net_1 ), .Y(data_buf6_i_net_1));
    SLE \data_buf[0]  (.D(sound_card_ctrl_0), .CLK(sdclk_n_1), .EN(
        data_buf6_i_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_buf[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  update_strobe_RNO (.A(
        \update_ack_dly[1]_net_1 ), .Y(\update_ack_dly_i[1] ));
    SLE \update_ack_dly[1]  (.D(\update_ack_dly[0]_net_1 ), .CLK(
        sdclk_n_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[1]_net_1 ));
    SLE \update_strobe_dly[2]  (.D(\update_strobe_dly[1]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[2]_net_1 ));
    SLE \update_strobe_dly[0]  (.D(update_strobe_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[0]_net_1 ));
    SLE \update_strobe_dly[3]  (.D(\update_strobe_dly[2]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[3]_net_1 ));
    SLE \update_ack_dly[0]  (.D(update_ack_net_1), .CLK(sdclk_n_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[0]_net_1 ));
    SLE update_ack (.D(\update_strobe_dly[3]_net_1 ), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        update_ack_net_1));
    CFG2 #( .INIT(4'h6) )  un1_update_strobe_dly (.A(update_ack_net_1), 
        .B(\update_strobe_dly[3]_net_1 ), .Y(un1_update_strobe_dly_0));
    SLE \update_strobe_dly[1]  (.D(\update_strobe_dly[0]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[1]_net_1 ));
    
endmodule


module sync_logic_3s(
       sound_card_ctrl,
       sdctrl_bck_divider,
       mclk_1,
       sdclk_n_1,
       N_4047_i
    );
input  [2:0] sound_card_ctrl;
output [2:0] sdctrl_bck_divider;
input  mclk_1;
input  sdclk_n_1;
input  N_4047_i;

    wire \update_ack_dly[1]_net_1 , \update_ack_dly_i[1] , 
        \update_ack_dly[0]_net_1 , VCC_net_1, update_ack_net_1, 
        GND_net_1, \update_strobe_dly[0]_net_1 , update_strobe_net_1, 
        \update_strobe_dly[1]_net_1 , \update_strobe_dly[2]_net_1 , 
        \update_strobe_dly[3]_net_1 , data_buf_sync_47_net_1, 
        data_buf_sync_48_net_1, data_buf_sync_49_net_1, 
        \data_buf[0]_net_1 , data_buf17_i_net_1, \data_buf[1]_net_1 , 
        \data_buf[2]_net_1 ;
    
    CFG1 #( .INIT(2'h1) )  update_strobe_RNO (.A(
        \update_ack_dly[1]_net_1 ), .Y(\update_ack_dly_i[1] ));
    SLE \data_buf[2]  (.D(sound_card_ctrl[2]), .CLK(sdclk_n_1), .EN(
        data_buf17_i_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_buf[2]_net_1 ));
    SLE \data_buf[0]  (.D(sound_card_ctrl[0]), .CLK(sdclk_n_1), .EN(
        data_buf17_i_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_buf[0]_net_1 ));
    CFG4 #( .INIT(16'hCAAC) )  data_buf_sync_49 (.A(
        \data_buf[2]_net_1 ), .B(sdctrl_bck_divider[2]), .C(
        \update_strobe_dly[3]_net_1 ), .D(update_ack_net_1), .Y(
        data_buf_sync_49_net_1));
    SLE \update_ack_dly[0]  (.D(update_ack_net_1), .CLK(sdclk_n_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[0]_net_1 ));
    SLE \update_strobe_dly[3]  (.D(\update_strobe_dly[2]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[3]_net_1 ));
    SLE \update_strobe_dly[2]  (.D(\update_strobe_dly[1]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hCAAC) )  data_buf_sync_48 (.A(
        \data_buf[1]_net_1 ), .B(sdctrl_bck_divider[1]), .C(
        \update_strobe_dly[3]_net_1 ), .D(update_ack_net_1), .Y(
        data_buf_sync_48_net_1));
    SLE update_ack (.D(\update_strobe_dly[3]_net_1 ), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        update_ack_net_1));
    SLE \update_ack_dly[1]  (.D(\update_ack_dly[0]_net_1 ), .CLK(
        sdclk_n_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[1]_net_1 ));
    SLE \update_strobe_dly[1]  (.D(\update_strobe_dly[0]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[1]_net_1 ));
    SLE \data_buf_sync[0]  (.D(data_buf_sync_47_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdctrl_bck_divider[0]));
    SLE \data_buf_sync[1]  (.D(data_buf_sync_48_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdctrl_bck_divider[1]));
    VCC VCC (.Y(VCC_net_1));
    SLE \update_strobe_dly[0]  (.D(update_strobe_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[0]_net_1 ));
    CFG4 #( .INIT(16'hE4D8) )  data_buf_sync_47 (.A(
        \update_strobe_dly[3]_net_1 ), .B(\data_buf[0]_net_1 ), .C(
        sdctrl_bck_divider[0]), .D(update_ack_net_1), .Y(
        data_buf_sync_47_net_1));
    SLE \data_buf_sync[2]  (.D(data_buf_sync_49_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdctrl_bck_divider[2]));
    SLE \data_buf[1]  (.D(sound_card_ctrl[1]), .CLK(sdclk_n_1), .EN(
        data_buf17_i_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_buf[1]_net_1 ));
    SLE update_strobe (.D(\update_ack_dly_i[1] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(update_strobe_net_1));
    CFG2 #( .INIT(4'h9) )  data_buf17_i (.A(update_strobe_net_1), .B(
        \update_ack_dly[1]_net_1 ), .Y(data_buf17_i_net_1));
    
endmodule


module bigfifo(
       test_0_HADDR,
       test_0_HWDATA,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0,
       dout,
       status,
       din,
       bus_state_0,
       state_0_0,
       state_0_d0,
       test_0_HTRANS_0,
       test_0_HADDR_i_0,
       buffer_under_runlde_0_a6_2,
       wen,
       read_en,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       test_0_HWRITE,
       sdclk_n_1,
       is_last_data,
       N_4047_i,
       mclk_1
    );
output [16:2] test_0_HADDR;
output [31:0] test_0_HWDATA;
input  [31:0] u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0;
output [31:0] dout;
output [7:6] status;
input  [31:0] din;
input  bus_state_0;
input  state_0_0;
input  state_0_d0;
output test_0_HTRANS_0;
output test_0_HADDR_i_0;
output buffer_under_runlde_0_a6_2;
input  wen;
input  read_en;
input  u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
output test_0_HWRITE;
input  sdclk_n_1;
input  is_last_data;
input  N_4047_i;
input  mclk_1;

    wire fifo_level, \write_addr_i[0] , \c1[26]_net_1 , VCC_net_1, 
        \c0[26]_net_1 , GND_net_1, \c1[27]_net_1 , \c0[27]_net_1 , 
        \c1[28]_net_1 , \c0[28]_net_1 , \c1[29]_net_1 , \c0[29]_net_1 , 
        \c1[30]_net_1 , \c0[30]_net_1 , \c1[31]_net_1 , \c0[31]_net_1 , 
        \j[0]_net_1 , N_3471_i, \j[1]_net_1 , N_3470_i, \j[2]_net_1 , 
        N_3469_i, \j[3]_net_1 , N_3468_i, \c1[11]_net_1 , 
        \c0[11]_net_1 , \c1[12]_net_1 , \c0[12]_net_1 , \c1[13]_net_1 , 
        \c0[13]_net_1 , \c1[14]_net_1 , \c0[14]_net_1 , \c1[15]_net_1 , 
        \c0[15]_net_1 , \c1[16]_net_1 , \c0[16]_net_1 , \c1[17]_net_1 , 
        \c0[17]_net_1 , \c1[18]_net_1 , \c0[18]_net_1 , \c1[19]_net_1 , 
        \c0[19]_net_1 , \c1[20]_net_1 , \c0[20]_net_1 , \c1[21]_net_1 , 
        \c0[21]_net_1 , \c1[22]_net_1 , \c0[22]_net_1 , \c1[23]_net_1 , 
        \c0[23]_net_1 , \c1[24]_net_1 , \c0[24]_net_1 , \c1[25]_net_1 , 
        \c0[25]_net_1 , \isl[0]_net_1 , \isl[1]_net_1 , \c1[0]_net_1 , 
        \c0[0]_net_1 , \c1[1]_net_1 , \c0[1]_net_1 , \c1[2]_net_1 , 
        \c0[2]_net_1 , \c1[3]_net_1 , \c0[3]_net_1 , \c1[4]_net_1 , 
        \c0[4]_net_1 , \c1[5]_net_1 , \c0[5]_net_1 , \c1[6]_net_1 , 
        \c0[6]_net_1 , \c1[7]_net_1 , \c0[7]_net_1 , \c1[8]_net_1 , 
        \c0[8]_net_1 , \c1[9]_net_1 , \c0[9]_net_1 , \c1[10]_net_1 , 
        \c0[10]_net_1 , N_3847_i, \a_full[0]_net_1 , full, 
        \a_full[1]_net_1 , \a_full[2]_net_1 , \a_empty[0]_net_1 , 
        empty_net_1, \a_empty[1]_net_1 , \a_empty[2]_net_1 , 
        \sync_wen[0]_net_1 , wen_toggle_net_1, \sync_wen[1]_net_1 , 
        \sync_wen[2]_net_1 , \n_HWDATA[30]_net_1 , un25_0_0_net_1, 
        \n_HWDATA[31]_net_1 , \n_HWDATA[15]_net_1 , 
        \n_HWDATA[16]_net_1 , \n_HWDATA[17]_net_1 , 
        \n_HWDATA[18]_net_1 , \n_HWDATA[19]_net_1 , 
        \n_HWDATA[20]_net_1 , \n_HWDATA[21]_net_1 , 
        \n_HWDATA[22]_net_1 , \n_HWDATA[23]_net_1 , 
        \n_HWDATA[24]_net_1 , \n_HWDATA[25]_net_1 , 
        \n_HWDATA[26]_net_1 , \n_HWDATA[27]_net_1 , 
        \n_HWDATA[28]_net_1 , \n_HWDATA[29]_net_1 , 
        \n_HWDATA[0]_net_1 , \n_HWDATA[1]_net_1 , \n_HWDATA[2]_net_1 , 
        \n_HWDATA[3]_net_1 , \n_HWDATA[4]_net_1 , \n_HWDATA[5]_net_1 , 
        \n_HWDATA[6]_net_1 , \n_HWDATA[7]_net_1 , \n_HWDATA[8]_net_1 , 
        \n_HWDATA[9]_net_1 , \n_HWDATA[10]_net_1 , 
        \n_HWDATA[11]_net_1 , \n_HWDATA[12]_net_1 , 
        \n_HWDATA[13]_net_1 , \n_HWDATA[14]_net_1 , 
        \read_addr[13]_net_1 , \read_addroi[13] , N_3845_i, 
        \addr[0]_net_1 , \n_addr[0] , N_272_i, \addr[1]_net_1 , 
        \n_addr[1] , \addr[2]_net_1 , \n_addr[2] , \addr[3]_net_1 , 
        \n_addr[3] , \addr[4]_net_1 , \n_addr[4] , \addr[5]_net_1 , 
        \n_addr[5] , \addr[6]_net_1 , \n_addr[6] , \addr[7]_net_1 , 
        \n_addr[7] , \addr[8]_net_1 , \n_addr[8] , \addr[9]_net_1 , 
        \n_addr[9] , \addr[10]_net_1 , \n_addr[10] , \addr[11]_net_1 , 
        \n_addr[11] , \addr[12]_net_1 , \n_addr[12] , \addr[13]_net_1 , 
        \n_addr[13] , \write_addr[12]_net_1 , \next_write_addr[12] , 
        N_126, \write_addr[13]_net_1 , \next_write_addr[13] , 
        \read_addr[0]_net_1 , read_addr_inc_s_1_419_Y, 
        \read_addr[1]_net_1 , \read_addroi[1] , \read_addr[2]_net_1 , 
        \read_addroi[2] , \read_addr[3]_net_1 , \read_addroi[3] , 
        \read_addr[4]_net_1 , \read_addroi[4] , \read_addr[5]_net_1 , 
        \read_addroi[5] , \read_addr[6]_net_1 , \read_addroi[6] , 
        \read_addr[7]_net_1 , \read_addroi[7] , \read_addr[8]_net_1 , 
        \read_addroi[8] , \read_addr[9]_net_1 , \read_addroi[9] , 
        \read_addr[10]_net_1 , \read_addroi[10] , 
        \read_addr[11]_net_1 , \read_addroi[11] , 
        \read_addr[12]_net_1 , \read_addroi[12] , 
        \write_block_addr[11]_net_1 , \next_write_addr[11] , 
        n_write_block_addr_0_sqmuxa, \write_block_addr[12]_net_1 , 
        \write_block_addr[13]_net_1 , \write_addr[1]_net_1 , 
        \next_write_addr[1] , \write_addr[2]_net_1 , 
        \next_write_addr[2] , \write_addr[3]_net_1 , 
        \next_write_addr[3] , \write_addr[4]_net_1 , 
        \next_write_addr[4] , \write_addr[5]_net_1 , 
        \next_write_addr[5] , \write_addr[6]_net_1 , 
        \next_write_addr[6] , \write_addr[7]_net_1 , 
        \next_write_addr[7] , \write_addr[8]_net_1 , 
        \next_write_addr[8] , \write_addr[9]_net_1 , 
        \next_write_addr[9] , \write_addr[10]_net_1 , 
        \next_write_addr[10] , \write_addr[11]_net_1 , 
        \write_block_addr[0]_net_1 , \write_block_addr[1]_net_1 , 
        \write_block_addr[2]_net_1 , \write_block_addr[3]_net_1 , 
        \write_block_addr[4]_net_1 , \write_block_addr[5]_net_1 , 
        \write_block_addr[6]_net_1 , \write_block_addr[7]_net_1 , 
        \write_block_addr[8]_net_1 , \write_block_addr[9]_net_1 , 
        \write_block_addr[10]_net_1 , N_729_i, un1_n_HWRITE_0_sqmuxa_3, 
        N_155_i_0_i, N_3846_i, un1_n_HWRITE_0_sqmuxa_4, N_274_i, 
        ready_net_1, \state[1]_net_1 , \state_ns[1] , \state[2]_net_1 , 
        \state_ns[2] , \state[3]_net_1 , \state[4]_net_1 , 
        \state_ns[4] , empty_2, \state[0]_net_1 , N_155_i_0, 
        wen_toggle_2_net_1, \i[0]_net_1 , \i_lm[0] , ie, \i[1]_net_1 , 
        \i_lm[1] , \i[2]_net_1 , \i_lm[2] , \i[3]_net_1 , \i_lm[3] , 
        \i[4]_net_1 , \i_lm[4] , \i[5]_net_1 , \i_lm[5] , \i[6]_net_1 , 
        \i_lm[6] , \i[7]_net_1 , \i_lm[7] , N_36_mux_reto, N_36_mux, 
        \fifo_level_reto[12] , \fifo_level[12] , \fifo_level_reto[13] , 
        \fifo_level[13] , \read_addr_inc_reti[13] , 
        \read_addr_inc_reti[12] , \read_addr_inc_reti[11] , 
        \read_addr_inc_reti[10] , \read_addr_inc_reti[9] , 
        \read_addr_inc_reti[8] , \read_addr_inc_reti[7] , 
        \read_addr_inc_reti[6] , \read_addr_inc_reti[5] , 
        \read_addr_inc_reti[4] , \read_addr_inc_reti[3] , 
        \read_addr_inc_reti[2] , \read_addr_inc_reti[1] , 
        fifo_level_cry_0_net_1, fifo_level_cry_0_Y, 
        fifo_level_cry_1_net_1, \fifo_level[1] , 
        fifo_level_cry_2_net_1, \fifo_level[2] , 
        fifo_level_cry_3_net_1, \fifo_level[3] , 
        fifo_level_cry_4_net_1, \fifo_level[4] , 
        fifo_level_cry_5_net_1, full_2lto5, fifo_level_cry_6_net_1, 
        \fifo_level[6] , fifo_level_cry_7_net_1, \fifo_level[7] , 
        fifo_level_cry_8_net_1, \fifo_level[8] , 
        fifo_level_cry_9_net_1, \fifo_level[9] , 
        fifo_level_cry_10_net_1, \fifo_level[10] , 
        fifo_level_cry_11_net_1, full_2lto11, fifo_level_cry_12_net_1, 
        \next_read_addr_0_data_tmp[0] , \next_read_addr_0_data_tmp[1] , 
        \next_read_addr_0_data_tmp[2] , \next_read_addr_0_data_tmp[3] , 
        \next_read_addr_0_data_tmp[4] , \next_read_addr_0_data_tmp[5] , 
        \next_read_addr_0_data_tmp[6] , i_s_416_FCO, \i_cry[1]_net_1 , 
        \i_s[1] , \i_cry[2]_net_1 , \i_s[2] , \i_cry[3]_net_1 , 
        \i_s[3] , \i_cry[4]_net_1 , \i_s[4] , \i_cry[5]_net_1 , 
        \i_s[5] , \i_s[7]_net_1 , \i_cry[6]_net_1 , \i_s[6] , 
        read_addr_inc_s_1_419_FCO, read_addr_inc_cry_1_net_1, 
        read_addr_inc_cry_2_net_1, read_addr_inc_cry_3_net_1, 
        read_addr_inc_cry_4_net_1, read_addr_inc_cry_5_net_1, 
        read_addr_inc_cry_6_net_1, read_addr_inc_cry_7_net_1, 
        read_addr_inc_cry_8_net_1, read_addr_inc_cry_9_net_1, 
        read_addr_inc_cry_10_net_1, read_addr_inc_cry_11_net_1, 
        read_addr_inc_cry_12_net_1, next_write_addr_s_1_420_FCO, 
        next_write_addr_cry_1_net_1, next_write_addr_cry_2_net_1, 
        next_write_addr_cry_3_net_1, next_write_addr_cry_4_net_1, 
        next_write_addr_cry_5_net_1, next_write_addr_cry_6_net_1, 
        next_write_addr_cry_7_net_1, next_write_addr_cry_8_net_1, 
        next_write_addr_cry_9_net_1, next_write_addr_cry_10_net_1, 
        next_write_addr_cry_11_net_1, next_write_addr_cry_12_net_1, 
        N_3489, n_d04_i_4_net_1, N_3484, N_3907, 
        n_d04_i_a3_RNI8AAV_net_1, N_3850, N_3886, N_3891, 
        un1_n_HWRITE_0_sqmuxa_7_0_2_net_1, n_d04_i_RNIVD122_net_1, 
        n_d04_i_4_N_2L1_net_1, n_d04_i_4_N_3L3_net_1, 
        n_d04_i_4_N_4L5_net_1, N_3474, 
        un1_n_HWRITE_0_sqmuxa_7_0_2_1_net_1, N_25_mux, m20_1, 
        fifo_level_cry_5_RNI5KEJ_net_1, 
        fifo_level_cry_10_RNIIKKL1_net_1, m13_5, m13_1, N_285_i, 
        \n_addr_iv_0_a2_0[13]_net_1 , m20_e_1, 
        un1_state_2_0_a2_2_6_a3_3_net_1, \state_ns_0_a3_0_1[1]_net_1 , 
        N_3472, N_3478, N_3888, N_3853, N_246_i, 
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_0_2, 
        un1_state_2_0_a2_2_6_a3_4_net_1, N_3475, N_3482, ilde_0_1, 
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_1_0, N_3477, N_3849, 
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_0_4, 
        un1_n_HWRITE_1_sqmuxa_2_i_0_233_i_o3_i_o2_d, N_3467, 
        un1_state_5;
    
    SLE \c0[22]  (.D(din[22]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[22]_net_1 ));
    CFG2 #( .INIT(4'h6) )  wen_toggle_2 (.A(wen_toggle_net_1), .B(wen), 
        .Y(wen_toggle_2_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[10]  (.A(
        \write_addr[10]_net_1 ), .B(\read_addr[10]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[10] ));
    SLE \state[0]  (.D(N_155_i_0), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    SLE \c0[24]  (.D(din[24]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[24]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[3]  (.A(\addr[1]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[3]));
    SLE \d0[9]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[9]));
    CFG2 #( .INIT(4'hE) )  \HADDR_2[7]  (.A(\addr[5]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[7]));
    SLE \addr[11]  (.D(\n_addr[11] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[11]_net_1 ));
    SLE \i[7]  (.D(\i_lm[7] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[7]_net_1 ));
    SLE \HWDATA[5]  (.D(\n_HWDATA[5]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[5]));
    SLE \c0[6]  (.D(din[6]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[6]_net_1 ));
    SLE \addr[7]  (.D(\n_addr[7] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[7]_net_1 ));
    SLE \d0[25]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[25]));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_10 (.A(VCC_net_1), 
        .B(\write_addr[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_9_net_1), .S(\next_write_addr[10] ), .Y(), 
        .FCO(next_write_addr_cry_10_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[0]  (.A(\state[2]_net_1 ), 
        .B(N_3849), .C(\read_addr[0]_net_1 ), .D(fifo_level), .Y(
        \n_addr[0] ));
    SLE \c1[3]  (.D(\c0[3]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[3]_net_1 ));
    SLE \c1[13]  (.D(\c0[13]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[13]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  un1_state_2_0_a2_2_6_a3 (.A(
        \i[5]_net_1 ), .B(\i[7]_net_1 ), .C(
        un1_state_2_0_a2_2_6_a3_4_net_1), .D(
        un1_state_2_0_a2_2_6_a3_3_net_1), .Y(N_285_i));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_8 (.A(VCC_net_1), 
        .B(\write_addr[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_7_net_1), .S(\next_write_addr[8] ), .Y(), 
        .FCO(next_write_addr_cry_8_net_1));
    CFG4 #( .INIT(16'hFBAA) )  \n_addr_iv_0_o2[13]  (.A(
        \state[1]_net_1 ), .B(\state[0]_net_1 ), .C(N_285_i), .D(
        \n_addr_iv_0_a2_0[13]_net_1 ), .Y(N_3849));
    SLE \write_addr[2]  (.D(\next_write_addr[2] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[2]_net_1 ));
    SLE \d0[5]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_12 (.A(VCC_net_1), 
        .B(\read_addroi[12] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_11_net_1), .S(\read_addr_inc_reti[12] ), .Y()
        , .FCO(read_addr_inc_cry_12_net_1));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_10 (.A(VCC_net_1), 
        .B(\read_addroi[10] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_9_net_1), .S(\read_addr_inc_reti[10] ), .Y(), 
        .FCO(read_addr_inc_cry_10_net_1));
    CFG2 #( .INIT(4'h8) )  pipeline_cmd_RNO (.A(N_285_i), .B(
        \state[0]_net_1 ), .Y(N_729_i));
    SLE \i[0]  (.D(\i_lm[0] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[0]_net_1 ));
    SLE \d0[1]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[1]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[14]  (.A(\state[0]_net_1 ), .B(
        \c1[14]_net_1 ), .Y(\n_HWDATA[14]_net_1 ));
    ARI1 #( .INIT(20'h68421) )  \write_block_addr_RNIFCED3[6]  (.A(
        \write_block_addr[7]_net_1 ), .B(\read_addroi[6] ), .C(
        \read_addroi[7] ), .D(\write_block_addr[6]_net_1 ), .FCI(
        \next_read_addr_0_data_tmp[2] ), .S(), .Y(), .FCO(
        \next_read_addr_0_data_tmp[3] ));
    ARI1 #( .INIT(20'h68421) )  \write_block_addr_RNI38V31[2]  (.A(
        \write_block_addr[3]_net_1 ), .B(\read_addroi[2] ), .C(
        \read_addroi[3] ), .D(\write_block_addr[2]_net_1 ), .FCI(
        \next_read_addr_0_data_tmp[0] ), .S(), .Y(), .FCO(
        \next_read_addr_0_data_tmp[1] ));
    SLE \d0[19]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[19]));
    CFG2 #( .INIT(4'h1) )  un1_state_2_0_a2_2_6_a3_3 (.A(\i[4]_net_1 ), 
        .B(\i[3]_net_1 ), .Y(un1_state_2_0_a2_2_6_a3_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_5 (.A(VCC_net_1), .B(
        \read_addroi[5] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_4_net_1), .S(\read_addr_inc_reti[5] ), .Y(), 
        .FCO(read_addr_inc_cry_5_net_1));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_5 (.A(
        \write_addr[5]_net_1 ), .B(\read_addr[5]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_4_net_1), .S(full_2lto5), 
        .Y(), .FCO(fifo_level_cry_5_net_1));
    SLE \c0[13]  (.D(din[13]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[13]_net_1 ));
    SLE \write_addr[0]  (.D(\write_addr_i[0] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(fifo_level));
    SLE \read_addr[1]  (.D(\read_addroi[1] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[1]_net_1 ));
    SLE \d0[24]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[24]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[19]  (.A(\state[0]_net_1 ), .B(
        \c1[19]_net_1 ), .Y(\n_HWDATA[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_9 (.A(VCC_net_1), .B(
        \read_addroi[9] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_8_net_1), .S(\read_addr_inc_reti[9] ), .Y(), 
        .FCO(read_addr_inc_cry_9_net_1));
    SLE \c1[19]  (.D(\c0[19]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[19]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[10]  (.A(\addr[8]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[10]));
    CFG4 #( .INIT(16'hAA03) )  \i_lm_0[2]  (.A(\i_s[2] ), .B(N_3891), 
        .C(un1_n_HWRITE_0_sqmuxa_7_0_2_net_1), .D(
        n_d04_i_RNIVD122_net_1), .Y(\i_lm[2] ));
    SLE \HWDATA[2]  (.D(\n_HWDATA[2]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[2]));
    CFG4 #( .INIT(16'h2F00) )  fifo_level_cry_0_RNITJKL1 (.A(
        fifo_level_cry_0_Y), .B(\fifo_level[1] ), .C(\fifo_level[2] ), 
        .D(fifo_level_cry_5_RNI5KEJ_net_1), .Y(N_25_mux));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_4 (.A(VCC_net_1), 
        .B(\write_addr[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_3_net_1), .S(\next_write_addr[4] ), .Y(), 
        .FCO(next_write_addr_cry_4_net_1));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[6]  (.A(\state[0]_net_1 ), .B(
        \c1[6]_net_1 ), .Y(\n_HWDATA[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_8 (.A(VCC_net_1), .B(
        \read_addroi[8] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_7_net_1), .S(\read_addr_inc_reti[8] ), .Y(), 
        .FCO(read_addr_inc_cry_8_net_1));
    SLE \d0[13]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[13]));
    SLE \c1[26]  (.D(\c0[26]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[26]_net_1 ));
    SLE \c0[19]  (.D(din[19]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[19]_net_1 ));
    SLE \d0[22]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[22]));
    CFG2 #( .INIT(4'hE) )  un1_state_4_0_i_o2 (.A(\state[2]_net_1 ), 
        .B(\state[3]_net_1 ), .Y(N_3850));
    SLE \d0[17]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[17]));
    SLE \sync_wen[2]  (.D(\sync_wen[1]_net_1 ), .CLK(mclk_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\sync_wen[2]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \n_j_i_o3_0[1]  (.A(\j[2]_net_1 ), .B(
        \j[3]_net_1 ), .Y(N_3478));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[13]  (.A(
        \write_addr[13]_net_1 ), .B(\read_addr[13]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[13] ));
    CFG4 #( .INIT(16'h00FE) )  \state_RNI88781[3]  (.A(
        \state[1]_net_1 ), .B(\state[2]_net_1 ), .C(\state[3]_net_1 ), 
        .D(read_en), .Y(un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_1_0));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[5]  (.A(
        \write_addr[5]_net_1 ), .B(\read_addr[5]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[5] ));
    SLE \c0[9]  (.D(din[9]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[9]_net_1 ));
    SLE read_addr_ret_2 (.D(\read_addr_inc_reti[11] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[11] ));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[8]  (.A(
        \write_addr[8]_net_1 ), .B(\read_addr[8]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[8] ));
    SLE \HWDATA[3]  (.D(\n_HWDATA[3]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[3]));
    SLE \d0[18]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[18]));
    SLE \a_empty[3]  (.D(\a_empty[2]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(status[6]));
    SLE \j[3]  (.D(N_3468_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\j[3]_net_1 ));
    SLE \write_addr[11]  (.D(\next_write_addr[11] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[11]_net_1 ));
    SLE \state[4]  (.D(\state_ns[4] ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[4]_net_1 ));
    SLE \c1[6]  (.D(\c0[6]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[6]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \HADDR_2[15]  (.A(\addr[13]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[15]));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_0 (.A(fifo_level), .B(
        \read_addr[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(fifo_level_cry_0_Y), .FCO(
        fifo_level_cry_0_net_1));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[27]  (.A(\state[0]_net_1 ), .B(
        \c1[27]_net_1 ), .Y(\n_HWDATA[27]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[20]  (.A(\state[0]_net_1 ), .B(
        \c1[20]_net_1 ), .Y(\n_HWDATA[20]_net_1 ));
    SLE read_addr_ret_4 (.D(\read_addr_inc_reti[9] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[9] ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_7 (.A(VCC_net_1), .B(
        \read_addroi[7] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_6_net_1), .S(\read_addr_inc_reti[7] ), .Y(), 
        .FCO(read_addr_inc_cry_7_net_1));
    CFG3 #( .INIT(8'h51) )  \HTRANS_1_RNO[1]  (.A(\state[4]_net_1 ), 
        .B(N_3850), .C(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .Y(
        N_3846_i));
    SLE \d0[26]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[26]));
    SLE \read_addr[7]  (.D(\read_addroi[7] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[7]_net_1 ));
    SLE \c1[21]  (.D(\c0[21]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[21]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[3]  (.A(\state[0]_net_1 ), .B(
        \c1[3]_net_1 ), .Y(\n_HWDATA[3]_net_1 ));
    SLE \c1[15]  (.D(\c0[15]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[15]_net_1 ));
    SLE \addr[0]  (.D(\n_addr[0] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[0]_net_1 ));
    CFG4 #( .INIT(16'hC844) )  \j_RNO[2]  (.A(N_3475), .B(un1_state_5), 
        .C(\j[3]_net_1 ), .D(\j[2]_net_1 ), .Y(N_3469_i));
    SLE \c0[5]  (.D(din[5]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[5]_net_1 ));
    SLE read_addr_ret_7 (.D(\read_addr_inc_reti[6] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[6] ));
    SLE \HWDATA[17]  (.D(\n_HWDATA[17]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[17]));
    SLE \c1[2]  (.D(\c0[2]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[2]_net_1 ));
    SLE \write_addr[13]  (.D(\next_write_addr[13] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[13]_net_1 ));
    SLE \c1[10]  (.D(\c0[10]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[10]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[13]  (.A(\state[0]_net_1 ), .B(
        \c1[13]_net_1 ), .Y(\n_HWDATA[13]_net_1 ));
    SLE \c0[1]  (.D(din[1]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[1]_net_1 ));
    SLE \a_full[3]  (.D(\a_full[2]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(status[7]));
    SLE \d0[2]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[2]));
    SLE \addr[8]  (.D(\n_addr[8] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[8]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \state_ns_0_a3_0_1[1]  (.A(\state[2]_net_1 )
        , .B(\state[0]_net_1 ), .Y(\state_ns_0_a3_0_1[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_3 (.A(VCC_net_1), .B(
        \read_addroi[3] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_2_net_1), .S(\read_addr_inc_reti[3] ), .Y(), 
        .FCO(read_addr_inc_cry_3_net_1));
    SLE \c0[31]  (.D(din[31]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[31]_net_1 ));
    SLE \c0[15]  (.D(din[15]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[15]_net_1 ));
    SLE pipeline_cmd (.D(N_729_i), .CLK(mclk_1), .EN(
        un1_n_HWRITE_0_sqmuxa_3), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HADDR[16]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[28]  (.A(\state[0]_net_1 ), .B(
        \c1[28]_net_1 ), .Y(\n_HWDATA[28]_net_1 ));
    SLE \d0[11]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[11]));
    SLE \write_block_addr[3]  (.D(\next_write_addr[3] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[3]_net_1 ));
    CFG2 #( .INIT(4'hB) )  \n_j_i_o3[0]  (.A(N_3478), .B(\j[1]_net_1 ), 
        .Y(N_3482));
    CFG3 #( .INIT(8'h70) )  \state_ns_i_o2_i_a3[0]  (.A(N_285_i), .B(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .C(\state[0]_net_1 )
        , .Y(N_155_i_0));
    SLE \d0[20]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[20]));
    SLE read_addr_ret_6 (.D(\read_addr_inc_reti[7] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[7] ));
    SLE \c0[10]  (.D(din[10]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[10]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[2]  (.A(
        \write_addr[2]_net_1 ), .B(\read_addr[2]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[2] ));
    SLE \c1[18]  (.D(\c0[18]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[18]_net_1 ));
    SLE \write_addr[3]  (.D(\next_write_addr[3] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[3]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[1]  (.A(
        \write_addr[1]_net_1 ), .B(\read_addr[1]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[1] ));
    SLE ready (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .CLK(
        mclk_1), .EN(\state[1]_net_1 ), .ALn(N_4047_i), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        ready_net_1));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[14]  (.A(\addr[12]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[14]));
    SLE read_addr_ret_11 (.D(\read_addr_inc_reti[2] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[2] ));
    SLE \c0[27]  (.D(din[27]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[27]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[22]  (.A(\state[0]_net_1 ), .B(
        \c1[22]_net_1 ), .Y(\n_HWDATA[22]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[9]  (.A(\addr[7]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[9]));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_4 (.A(
        \write_addr[4]_net_1 ), .B(\read_addr[4]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_3_net_1), .S(
        \fifo_level[4] ), .Y(), .FCO(fifo_level_cry_4_net_1));
    SLE \c1[23]  (.D(\c0[23]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[23]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[21]  (.A(\state[0]_net_1 ), .B(
        \c1[21]_net_1 ), .Y(\n_HWDATA[21]_net_1 ));
    SLE \c0[18]  (.D(din[18]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[18]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[12]  (.A(
        \write_addr[12]_net_1 ), .B(\read_addr[12]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[12] ));
    SLE \write_block_addr[6]  (.D(\next_write_addr[6] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[6]_net_1 ));
    SLE \write_block_addr[5]  (.D(\next_write_addr[5] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[5]_net_1 ));
    SLE \write_block_addr[11]  (.D(\next_write_addr[11] ), .CLK(mclk_1)
        , .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[11]_net_1 ));
    SLE \HWDATA[27]  (.D(\n_HWDATA[27]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[27]));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[11]  (.A(\addr[9]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[11]));
    SLE \addr[5]  (.D(\n_addr[5] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[5]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \HWDATA[8]  (.D(\n_HWDATA[8]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[8]));
    SLE \read_addr[13]  (.D(\read_addroi[13] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[13]_net_1 ));
    CFG4 #( .INIT(16'h004C) )  n_d04_i_4_RNIGKLK1 (.A(n_d04_i_4_net_1), 
        .B(n_d04_i_a3_RNI8AAV_net_1), .C(\state[1]_net_1 ), .D(N_3850), 
        .Y(N_3886));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[6]  (.A(\addr[4]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[6]));
    CFG2 #( .INIT(4'hE) )  un1_n_HWRITE_0_sqmuxa_4_0_1 (.A(N_3891), .B(
        N_126), .Y(un1_n_HWRITE_0_sqmuxa_4));
    SLE \sync_wen[1]  (.D(\sync_wen[0]_net_1 ), .CLK(mclk_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\sync_wen[1]_net_1 ));
    SLE \HWDATA[18]  (.D(\n_HWDATA[18]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[18]));
    SLE \c1[29]  (.D(\c0[29]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[29]_net_1 ));
    SLE \write_addr[6]  (.D(\next_write_addr[6] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[6]_net_1 ));
    SLE \write_addr[5]  (.D(\next_write_addr[5] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[5]_net_1 ));
    SLE \read_addr[12]  (.D(\read_addroi[12] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  i_s_416 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(i_s_416_FCO));
    SLE \addr[1]  (.D(\n_addr[1] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[1]_net_1 ));
    SLE \d0[0]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[0]));
    SLE \read_addr[5]  (.D(\read_addroi[5] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[12]  (.A(\addr[10]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[12]));
    CFG4 #( .INIT(16'hC080) )  un1_state_4_0_i_o2_RNIBB713 (.A(
        \state[1]_net_1 ), .B(
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_0_2), .C(N_3477), .D(
        N_3850), .Y(un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_0_4));
    CFG3 #( .INIT(8'h8F) )  \state_ns_i_o2_i_a3_i[0]  (.A(N_285_i), .B(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .C(\state[0]_net_1 )
        , .Y(N_155_i_0_i));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[8]  (.A(\addr[6]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[8]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[7]  (.A(\state[0]_net_1 ), .B(
        \c1[7]_net_1 ), .Y(\n_HWDATA[7]_net_1 ));
    SLE \HWDATA[15]  (.D(\n_HWDATA[15]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[15]));
    SLE read_addr_ret_12 (.D(\read_addr_inc_reti[1] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[1] ));
    CFG4 #( .INIT(16'h84C4) )  \j_RNO[1]  (.A(N_3472), .B(un1_state_5), 
        .C(\j[1]_net_1 ), .D(N_3478), .Y(N_3470_i));
    CFG2 #( .INIT(4'h1) )  fifo_level_cry_5_RNI5KEJ (.A(full_2lto11), 
        .B(full_2lto5), .Y(fifo_level_cry_5_RNI5KEJ_net_1));
    SLE \sync_wen[0]  (.D(wen_toggle_net_1), .CLK(mclk_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\sync_wen[0]_net_1 ));
    ARI1 #( .INIT(20'h49900) )  fifo_level_s_13 (.A(VCC_net_1), .B(
        \read_addr[13]_net_1 ), .C(\write_addr[13]_net_1 ), .D(
        GND_net_1), .FCI(fifo_level_cry_12_net_1), .S(\fifo_level[13] )
        , .Y(), .FCO());
    CFG2 #( .INIT(4'h7) )  \n_j_i_o3[1]  (.A(\state[1]_net_1 ), .B(
        \j[0]_net_1 ), .Y(N_3472));
    SLE \HWDATA[14]  (.D(\n_HWDATA[14]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[14]));
    SLE \write_addr[12]  (.D(\next_write_addr[12] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[12]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[5]  (.A(\state[0]_net_1 ), .B(
        \c1[5]_net_1 ), .Y(\n_HWDATA[5]_net_1 ));
    SLE \c0[2]  (.D(din[2]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[2]_net_1 ));
    SLE \write_block_addr[10]  (.D(\next_write_addr[10] ), .CLK(mclk_1)
        , .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[10]_net_1 ));
    SLE \c1[12]  (.D(\c0[12]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[12]_net_1 ));
    SLE \read_addr[8]  (.D(\read_addroi[8] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[8]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_3 (.A(
        \write_addr[3]_net_1 ), .B(\read_addr[3]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_2_net_1), .S(
        \fifo_level[3] ), .Y(), .FCO(fifo_level_cry_3_net_1));
    SLE \c1[14]  (.D(\c0[14]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[14]_net_1 ));
    SLE \write_block_addr[2]  (.D(\next_write_addr[2] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[2]_net_1 ));
    SLE \isl[1]  (.D(\isl[0]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\isl[1]_net_1 ));
    CFG4 #( .INIT(16'hE2CC) )  full_ret_RNO (.A(N_25_mux), .B(m20_1), 
        .C(fifo_level_cry_5_RNI5KEJ_net_1), .D(
        fifo_level_cry_10_RNIIKKL1_net_1), .Y(N_36_mux));
    ARI1 #( .INIT(20'h68421) )  \write_block_addr_RNIL46I4[8]  (.A(
        \write_block_addr[9]_net_1 ), .B(\read_addroi[8] ), .C(
        \read_addroi[9] ), .D(\write_block_addr[8]_net_1 ), .FCI(
        \next_read_addr_0_data_tmp[3] ), .S(), .Y(), .FCO(
        \next_read_addr_0_data_tmp[4] ));
    SLE \c1[5]  (.D(\c0[5]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[5]_net_1 ));
    SLE read_addr_ret_10 (.D(\read_addr_inc_reti[3] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[3] ));
    CFG4 #( .INIT(16'hB3A0) )  \state_ns_0[2]  (.A(\state[1]_net_1 ), 
        .B(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .C(N_246_i), .D(
        \state[2]_net_1 ), .Y(\state_ns[2] ));
    SLE read_addr_ret_1 (.D(\read_addr_inc_reti[12] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[12] ));
    SLE \HWDATA[4]  (.D(\n_HWDATA[4]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[4]));
    SLE \c0[12]  (.D(din[12]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_9 (.A(VCC_net_1), 
        .B(\write_addr[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_8_net_1), .S(\next_write_addr[9] ), .Y(), 
        .FCO(next_write_addr_cry_9_net_1));
    CFG2 #( .INIT(4'hB) )  \n_j_i_o3[2]  (.A(N_3472), .B(\j[1]_net_1 ), 
        .Y(N_3475));
    CFG4 #( .INIT(16'hE000) )  n_d04_i_a3 (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(\i[5]_net_1 ), .D(\i[4]_net_1 ), .Y(N_3484));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[9]  (.A(\state[0]_net_1 ), .B(
        \c1[9]_net_1 ), .Y(\n_HWDATA[9]_net_1 ));
    SLE \d0[7]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[7]));
    SLE \c0[14]  (.D(din[14]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[14]_net_1 ));
    SLE \HWDATA[7]  (.D(\n_HWDATA[7]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[7]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[24]  (.A(\state[0]_net_1 ), .B(
        \c1[24]_net_1 ), .Y(\n_HWDATA[24]_net_1 ));
    SLE \write_block_addr[4]  (.D(\next_write_addr[4] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[4]_net_1 ));
    SLE \c0[26]  (.D(din[26]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[26]_net_1 ));
    ARI1 #( .INIT(20'h68421) )  \write_block_addr_RNIEAU77[12]  (.A(
        \write_block_addr[13]_net_1 ), .B(\read_addroi[12] ), .C(
        \read_addroi[13] ), .D(\write_block_addr[12]_net_1 ), .FCI(
        \next_read_addr_0_data_tmp[5] ), .S(), .Y(), .FCO(
        \next_read_addr_0_data_tmp[6] ));
    CFG4 #( .INIT(16'h1000) )  \a_empty_RNIEFL71[3]  (.A(state_0_d0), 
        .B(state_0_0), .C(status[6]), .D(bus_state_0), .Y(
        buffer_under_runlde_0_a6_2));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[11]  (.A(
        \write_addr[11]_net_1 ), .B(\read_addr[11]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[11] ));
    SLE \HWDATA[0]  (.D(\n_HWDATA[0]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[0]));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[3]  (.A(n_d04_i_RNIVD122_net_1), .B(
        \i_s[3] ), .Y(\i_lm[3] ));
    SLE \HWDATA[28]  (.D(\n_HWDATA[28]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[28]));
    SLE \write_addr[10]  (.D(\next_write_addr[10] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[10]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_11 (.A(VCC_net_1), 
        .B(\read_addroi[11] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_10_net_1), .S(\read_addr_inc_reti[11] ), .Y()
        , .FCO(read_addr_inc_cry_11_net_1));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[29]  (.A(\state[0]_net_1 ), .B(
        \c1[29]_net_1 ), .Y(\n_HWDATA[29]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[0]  (.A(\state[0]_net_1 ), .B(
        \c1[0]_net_1 ), .Y(\n_HWDATA[0]_net_1 ));
    SLE \d0[15]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[15]));
    SLE \c1[25]  (.D(\c0[25]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[25]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_2 (.A(VCC_net_1), .B(
        \read_addroi[2] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_1_net_1), .S(\read_addr_inc_reti[2] ), .Y(), 
        .FCO(read_addr_inc_cry_2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_4 (.A(VCC_net_1), .B(
        \read_addroi[4] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_3_net_1), .S(\read_addr_inc_reti[4] ), .Y(), 
        .FCO(read_addr_inc_cry_4_net_1));
    SLE \HWDATA[11]  (.D(\n_HWDATA[11]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[11]));
    SLE \c1[31]  (.D(\c0[31]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[31]_net_1 ));
    SLE \HWDATA[25]  (.D(\n_HWDATA[25]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[25]));
    SLE \c1[20]  (.D(\c0[20]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[20]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_5 (.A(VCC_net_1), 
        .B(\write_addr[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_4_net_1), .S(\next_write_addr[5] ), .Y(), 
        .FCO(next_write_addr_cry_5_net_1));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_1 (.A(VCC_net_1), 
        .B(\write_addr[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_s_1_420_FCO), .S(\next_write_addr[1] ), .Y(), 
        .FCO(next_write_addr_cry_1_net_1));
    CFG4 #( .INIT(16'hF4FC) )  un1_state_2_0_a2_2_6_a3_RNI2RMB1 (.A(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .B(\state[0]_net_1 )
        , .C(N_3888), .D(N_285_i), .Y(ilde_0_1));
    SLE read_addr_ret_5 (.D(\read_addr_inc_reti[8] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[8] ));
    SLE \HWDATA[24]  (.D(\n_HWDATA[24]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[24]));
    CFG4 #( .INIT(16'h0004) )  n_d04_i_a3_RNIBTRQ (.A(N_3489), .B(
        \state[1]_net_1 ), .C(n_d04_i_4_net_1), .D(N_3484), .Y(
        N_3847_i));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[5]  (.A(\addr[3]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[5]));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[6]  (.A(n_d04_i_RNIVD122_net_1), .B(
        \i_s[6] ), .Y(\i_lm[6] ));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[2]  (.A(\addr[0]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[2]));
    SLE \addr[9]  (.D(\n_addr[9] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[9]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_6 (.A(VCC_net_1), .B(
        \read_addroi[6] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_5_net_1), .S(\read_addr_inc_reti[6] ), .Y(), 
        .FCO(read_addr_inc_cry_6_net_1));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_2 (.A(VCC_net_1), 
        .B(\write_addr[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_1_net_1), .S(\next_write_addr[2] ), .Y(), 
        .FCO(next_write_addr_cry_2_net_1));
    CFG2 #( .INIT(4'h8) )  fifo_level_cry_8_RNIVAPM (.A(
        \fifo_level[9] ), .B(\fifo_level[8] ), .Y(m20_e_1));
    SLE \d0[31]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[31]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[2]  (.A(\state[0]_net_1 ), .B(
        \c1[2]_net_1 ), .Y(\n_HWDATA[2]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  read_addr_inc_s_1_419 (.A(VCC_net_1), 
        .B(\read_addr[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(read_addr_inc_s_1_419_Y), .FCO(
        read_addr_inc_s_1_419_FCO));
    SLE \c0[0]  (.D(din[0]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_s[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[6]_net_1 ), .S(\i_s[7]_net_1 ), .Y(), .FCO());
    SLE \i[2]  (.D(\i_lm[2] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[2]_net_1 ));
    SLE \d0[8]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[8]));
    SLE \c0[21]  (.D(din[21]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[21]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_8 (.A(
        \write_addr[8]_net_1 ), .B(\read_addr[8]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_7_net_1), .S(
        \fifo_level[8] ), .Y(), .FCO(fifo_level_cry_8_net_1));
    SLE \c1[28]  (.D(\c0[28]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[28]_net_1 ));
    SLE \c0[30]  (.D(din[30]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[30]_net_1 ));
    SLE \d0[14]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[14]));
    CFG2 #( .INIT(4'hD) )  un1_state_5_0_o3_RNIER9I (.A(N_3853), .B(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .Y(N_272_i));
    SLE \HTRANS_1[1]  (.D(N_155_i_0_i), .CLK(mclk_1), .EN(N_3846_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(test_0_HTRANS_0));
    CFG1 #( .INIT(2'h1) )  \write_addr_RNITCFC[0]  (.A(fifo_level), .Y(
        \write_addr_i[0] ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[16]  (.A(\state[0]_net_1 ), .B(
        \c1[16]_net_1 ), .Y(\n_HWDATA[16]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[4]  (.A(\state[0]_net_1 ), .B(
        \c1[4]_net_1 ), .Y(\n_HWDATA[4]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  un1_n_HWRITE_0_sqmuxa_3_0_0 (.A(
        \state[4]_net_1 ), .B(N_3891), .C(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .Y(
        un1_n_HWRITE_0_sqmuxa_3));
    CFG3 #( .INIT(8'h01) )  n_read_addr_1_sqmuxa_i_a2 (.A(
        \state[1]_net_1 ), .B(\state[2]_net_1 ), .C(\state[3]_net_1 ), 
        .Y(N_3907));
    CFG4 #( .INIT(16'hAA03) )  \i_lm_0[1]  (.A(\i_s[1] ), .B(N_3891), 
        .C(un1_n_HWRITE_0_sqmuxa_7_0_2_net_1), .D(
        n_d04_i_RNIVD122_net_1), .Y(\i_lm[1] ));
    CFG4 #( .INIT(16'h80AA) )  un1_n_HWRITE_0_sqmuxa_7_0_2 (.A(read_en)
        , .B(\state[1]_net_1 ), .C(n_d04_i_4_net_1), .D(
        un1_n_HWRITE_0_sqmuxa_7_0_2_1_net_1), .Y(
        un1_n_HWRITE_0_sqmuxa_7_0_2_net_1));
    CFG4 #( .INIT(16'hFFFE) )  n_d04_i_a3_RNIVVGL (.A(N_3484), .B(
        N_3489), .C(n_d04_i_4_net_1), .D(N_3850), .Y(
        un1_n_HWRITE_1_sqmuxa_2_i_0_233_i_o3_i_o2_d));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[6]  (.A(
        \write_addr[6]_net_1 ), .B(\read_addr[6]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[6] ));
    SLE \HWDATA[31]  (.D(\n_HWDATA[31]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[31]));
    CFG3 #( .INIT(8'h80) )  un1_n_HWRITE_0_sqmuxa_3_0_0_a3 (.A(N_285_i)
        , .B(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .C(
        \state[0]_net_1 ), .Y(N_3891));
    SLE \write_block_addr[12]  (.D(\next_write_addr[12] ), .CLK(mclk_1)
        , .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_s_1_420 (.A(VCC_net_1), 
        .B(fifo_level), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(next_write_addr_s_1_420_FCO));
    SLE \HWDATA[13]  (.D(\n_HWDATA[13]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[13]));
    SLE \state[3]  (.D(\state[2]_net_1 ), .CLK(mclk_1), .EN(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\state[3]_net_1 ));
    CFG4 #( .INIT(16'h4CC0) )  \j_RNO[0]  (.A(N_3482), .B(un1_state_5), 
        .C(\j[0]_net_1 ), .D(\state[1]_net_1 ), .Y(N_3471_i));
    CFG4 #( .INIT(16'h0307) )  un1_n_HWRITE_0_sqmuxa_7_0_2_1 (.A(
        N_3489), .B(\state[1]_net_1 ), .C(N_3850), .D(N_3484), .Y(
        un1_n_HWRITE_0_sqmuxa_7_0_2_1_net_1));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_7 (.A(
        \write_addr[7]_net_1 ), .B(\read_addr[7]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_6_net_1), .S(
        \fifo_level[7] ), .Y(), .FCO(fifo_level_cry_7_net_1));
    SLE \d0[12]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[12]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[15]  (.A(\state[0]_net_1 ), .B(
        \c1[15]_net_1 ), .Y(\n_HWDATA[15]_net_1 ));
    ARI1 #( .INIT(20'h68421) )  \write_block_addr_RNI9OM82[4]  (.A(
        \write_block_addr[5]_net_1 ), .B(\read_addroi[4] ), .C(
        \read_addroi[5] ), .D(\write_block_addr[4]_net_1 ), .FCI(
        \next_read_addr_0_data_tmp[1] ), .S(), .Y(), .FCO(
        \next_read_addr_0_data_tmp[2] ));
    CFG3 #( .INIT(8'hFE) )  HWRITE_RNO (.A(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .B(\state[0]_net_1 )
        , .C(\state[1]_net_1 ), .Y(N_274_i));
    SLE \HWDATA[21]  (.D(\n_HWDATA[21]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[21]));
    SLE \i[6]  (.D(\i_lm[6] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(i_s_416_FCO), 
        .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    SLE \c0[7]  (.D(din[7]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[7]_net_1 ));
    CFG4 #( .INIT(16'h6444) )  \state_ns_0[4]  (.A(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .B(\state[4]_net_1 )
        , .C(N_3907), .D(N_285_i), .Y(\state_ns[4] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[4]  (.D(\i_lm[4] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[23]  (.A(\state[0]_net_1 ), .B(
        \c1[23]_net_1 ), .Y(\n_HWDATA[23]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un1_state_5_0_o3 (.A(\state[4]_net_1 ), .B(
        \state[3]_net_1 ), .Y(N_3853));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(\i_cry[6]_net_1 ));
    SLE \write_addr[1]  (.D(\next_write_addr[1] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[1]_net_1 ));
    SLE \HWDATA[16]  (.D(\n_HWDATA[16]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[16]));
    SLE \d0[29]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[29]));
    SLE \a_full[2]  (.D(\a_full[1]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\a_full[2]_net_1 ));
    SLE \d0[4]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[4]));
    SLE \c0[23]  (.D(din[23]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[23]_net_1 ));
    SLE read_addr_ret_8 (.D(\read_addr_inc_reti[5] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[5] ));
    CFG2 #( .INIT(4'h4) )  \n_addr_iv_0_a2_0[13]  (.A(\state[2]_net_1 )
        , .B(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .Y(
        \n_addr_iv_0_a2_0[13]_net_1 ));
    SLE \read_addr[6]  (.D(\read_addroi[6] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[6]_net_1 ));
    SLE \j[2]  (.D(N_3469_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\j[2]_net_1 ));
    SLE \write_addr[9]  (.D(\next_write_addr[9] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[9]_net_1 ));
    CFG3 #( .INIT(8'hDF) )  n_d04_i_o3_RNIN3DV (.A(\i[4]_net_1 ), .B(
        N_3474), .C(\i[3]_net_1 ), .Y(N_3477));
    SLE \d0[16]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[16]));
    SLE \a_full[1]  (.D(\a_full[0]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\a_full[1]_net_1 ));
    SLE \a_empty[1]  (.D(\a_empty[0]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\a_empty[1]_net_1 ));
    SLE \c1[9]  (.D(\c0[9]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[9]_net_1 ));
    SLE \c1[22]  (.D(\c0[22]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[22]_net_1 ));
    SLE \HWDATA[1]  (.D(\n_HWDATA[1]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[1]));
    SLE HWRITE (.D(un1_n_HWRITE_0_sqmuxa_4), .CLK(mclk_1), .EN(N_274_i)
        , .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(test_0_HWRITE));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[13]  (.A(\addr[11]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[13]));
    SLE \c1[24]  (.D(\c0[24]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[24]_net_1 ));
    CFG4 #( .INIT(16'hFF60) )  un25_0_0 (.A(\sync_wen[1]_net_1 ), .B(
        \sync_wen[2]_net_1 ), .C(\state[1]_net_1 ), .D(
        \state[0]_net_1 ), .Y(un25_0_0_net_1));
    CFG4 #( .INIT(16'hFF20) )  un1_state_5_0 (.A(\state[1]_net_1 ), .B(
        read_en), .C(N_3467), .D(N_3853), .Y(un1_state_5));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[3]  (.A(
        \write_addr[3]_net_1 ), .B(\read_addr[3]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[3] ));
    SLE \d0[23]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[23]));
    ARI1 #( .INIT(20'h64812) )  \write_block_addr_RNIFPLH[0]  (.A(
        \write_block_addr[1]_net_1 ), .B(\read_addr[0]_net_1 ), .C(
        \read_addroi[1] ), .D(\write_block_addr[0]_net_1 ), .FCI(
        GND_net_1), .S(), .Y(), .FCO(\next_read_addr_0_data_tmp[0] ));
    SLE \read_addr[3]  (.D(\read_addroi[3] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[3]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  un1_state_2_0_a2_2_6_a3_4 (.A(
        \i[6]_net_1 ), .B(\i[2]_net_1 ), .C(\i[1]_net_1 ), .D(
        \i[0]_net_1 ), .Y(un1_state_2_0_a2_2_6_a3_4_net_1));
    SLE \c0[29]  (.D(din[29]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[29]_net_1 ));
    SLE \write_addr[8]  (.D(\next_write_addr[8] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[8]_net_1 ));
    SLE \HWDATA[23]  (.D(\n_HWDATA[23]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[23]));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_6 (.A(
        \write_addr[6]_net_1 ), .B(\read_addr[6]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_5_net_1), .S(
        \fifo_level[6] ), .Y(), .FCO(fifo_level_cry_6_net_1));
    SLE \c1[8]  (.D(\c0[8]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[8]_net_1 ));
    SLE \c0[8]  (.D(din[8]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[8]_net_1 ));
    SLE \d0[27]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[27]));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[9]  (.A(
        \write_addr[9]_net_1 ), .B(\read_addr[9]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[9] ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_cry_1 (.A(VCC_net_1), .B(
        \read_addroi[1] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_s_1_419_FCO), .S(\read_addr_inc_reti[1] ), .Y(), 
        .FCO(read_addr_inc_cry_1_net_1));
    CFG4 #( .INIT(16'h2E0C) )  \state_ns_0[1]  (.A(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .B(\state[1]_net_1 )
        , .C(N_246_i), .D(\state_ns_0_a3_0_1[1]_net_1 ), .Y(
        \state_ns[1] ));
    CFG3 #( .INIT(8'h20) )  n_read_addr_1_sqmuxa_i_a2_RNI0NIN7 (.A(
        \next_read_addr_0_data_tmp[6] ), .B(N_3907), .C(read_en), .Y(
        N_3845_i));
    CFG4 #( .INIT(16'hFAF8) )  n_d04_i_RNIVD122 (.A(
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_1_0), .B(N_3850), .C(
        N_155_i_0), .D(N_3467), .Y(n_d04_i_RNIVD122_net_1));
    SLE \c1[1]  (.D(\c0[1]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[1]_net_1 ));
    SLE \c1[17]  (.D(\c0[17]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[17]_net_1 ));
    SLE empty (.D(empty_2), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(empty_net_1));
    CFG4 #( .INIT(16'hC4C0) )  \j_RNO[3]  (.A(N_3475), .B(un1_state_5), 
        .C(\j[3]_net_1 ), .D(\j[2]_net_1 ), .Y(N_3468_i));
    SLE \d0[10]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[10]));
    ARI1 #( .INIT(20'h68421) )  \write_block_addr_RNI97H06[10]  (.A(
        \write_block_addr[11]_net_1 ), .B(\read_addroi[10] ), .C(
        \read_addroi[11] ), .D(\write_block_addr[10]_net_1 ), .FCI(
        \next_read_addr_0_data_tmp[4] ), .S(), .Y(), .FCO(
        \next_read_addr_0_data_tmp[5] ));
    SLE read_addr_ret_9 (.D(\read_addr_inc_reti[4] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[4] ));
    CFG3 #( .INIT(8'h02) )  n_d04_i_4_N_3L3 (.A(ready_net_1), .B(
        \i[7]_net_1 ), .C(\i[6]_net_1 ), .Y(n_d04_i_4_N_3L3_net_1));
    SLE \d0[28]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[28]));
    SLE \addr[12]  (.D(\n_addr[12] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[12]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[7]  (.A(n_d04_i_RNIVD122_net_1), .B(
        \i_s[7]_net_1 ), .Y(\i_lm[7] ));
    SLE \d0[3]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[3]));
    SLE \addr[4]  (.D(\n_addr[4] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[4]_net_1 ));
    SLE \HWDATA[12]  (.D(\n_HWDATA[12]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[12]));
    SLE full_ret_2 (.D(\fifo_level[13] ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\fifo_level_reto[13] ));
    CFG4 #( .INIT(16'h8000) )  fifo_level_cry_10_RNIIKKL1 (.A(
        \fifo_level[6] ), .B(\fifo_level[7] ), .C(\fifo_level[10] ), 
        .D(m20_e_1), .Y(fifo_level_cry_10_RNIIKKL1_net_1));
    SLE \c1[0]  (.D(\c0[0]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[0]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \a_full_RNO[0]  (.A(\fifo_level_reto[13] ), 
        .B(\fifo_level_reto[12] ), .C(N_36_mux_reto), .Y(full));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    SLE \HWDATA[26]  (.D(\n_HWDATA[26]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[26]));
    SLE \addr[2]  (.D(\n_addr[2] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[2]_net_1 ));
    SLE \state[2]  (.D(\state_ns[2] ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_7 (.A(VCC_net_1), 
        .B(\write_addr[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_6_net_1), .S(\next_write_addr[7] ), .Y(), 
        .FCO(next_write_addr_cry_7_net_1));
    SLE \c0[17]  (.D(din[17]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[17]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_s_13 (.A(VCC_net_1), 
        .B(\write_addr[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_12_net_1), .S(\next_write_addr[13] ), .Y(), 
        .FCO());
    SLE \write_block_addr[1]  (.D(\next_write_addr[1] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[1]_net_1 ));
    SLE wen_toggle (.D(wen_toggle_2_net_1), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(wen_toggle_net_1));
    SLE \c1[4]  (.D(\c0[4]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[4]_net_1 ));
    SLE \read_addr[10]  (.D(\read_addroi[10] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[10]_net_1 ));
    SLE \addr[13]  (.D(\n_addr[13] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[13]_net_1 ));
    SLE \write_block_addr[7]  (.D(\next_write_addr[7] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[7]_net_1 ));
    SLE \isl[0]  (.D(is_last_data), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\isl[0]_net_1 ));
    SLE \addr[10]  (.D(\n_addr[10] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[10]_net_1 ));
    SLE \state[1]  (.D(\state_ns[1] ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[1]  (.A(\state[0]_net_1 ), .B(
        \c1[1]_net_1 ), .Y(\n_HWDATA[1]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  n_d04_i_o3 (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(\i[0]_net_1 ), .Y(N_3474));
    SLE \write_block_addr[9]  (.D(\next_write_addr[9] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[9]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[30]  (.A(\state[0]_net_1 ), .B(
        \c1[30]_net_1 ), .Y(\n_HWDATA[30]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_12 (.A(VCC_net_1), 
        .B(\write_addr[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_11_net_1), .S(\next_write_addr[12] ), .Y(), 
        .FCO(next_write_addr_cry_12_net_1));
    SLE \c1[30]  (.D(\c0[30]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[30]_net_1 ));
    SLE \i[5]  (.D(\i_lm[5] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[5]_net_1 ));
    CFG4 #( .INIT(16'h1115) )  n_d04_i_a3_RNI8AAV (.A(\state[4]_net_1 )
        , .B(\state[1]_net_1 ), .C(N_3489), .D(N_3484), .Y(
        n_d04_i_a3_RNI8AAV_net_1));
    CFG4 #( .INIT(16'h0001) )  \i_RNICPCI1[6]  (.A(\i[7]_net_1 ), .B(
        \i[6]_net_1 ), .C(\i[5]_net_1 ), .D(read_en), .Y(
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_0_2));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_2 (.A(
        \write_addr[2]_net_1 ), .B(\read_addr[2]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_1_net_1), .S(
        \fifo_level[2] ), .Y(), .FCO(fifo_level_cry_2_net_1));
    CFG4 #( .INIT(16'h0015) )  n_d04_i_4_N_2L1 (.A(\j[2]_net_1 ), .B(
        \j[1]_net_1 ), .C(\j[0]_net_1 ), .D(\j[3]_net_1 ), .Y(
        n_d04_i_4_N_2L1_net_1));
    SLE \write_block_addr[0]  (.D(\write_addr_i[0] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_11 (.A(VCC_net_1), 
        .B(\write_addr[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_10_net_1), .S(\next_write_addr[11] ), .Y(), 
        .FCO(next_write_addr_cry_11_net_1));
    SLE \c0[4]  (.D(din[4]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[4]_net_1 ));
    SLE \write_addr[4]  (.D(\next_write_addr[4] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[4]_net_1 ));
    SLE \HWDATA[10]  (.D(\n_HWDATA[10]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[10]));
    SLE \read_addr[11]  (.D(\read_addroi[11] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[11]_net_1 ));
    SLE \c0[25]  (.D(din[25]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[25]_net_1 ));
    SLE \HWDATA[19]  (.D(\n_HWDATA[19]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[19]));
    CFG4 #( .INIT(16'h2000) )  empty_RNO (.A(m13_5), .B(
        \fifo_level[13] ), .C(N_25_mux), .D(m13_1), .Y(empty_2));
    CFG4 #( .INIT(16'hAA03) )  \i_lm_0[5]  (.A(\i_s[5] ), .B(N_3891), 
        .C(un1_n_HWRITE_0_sqmuxa_7_0_2_net_1), .D(
        n_d04_i_RNIVD122_net_1), .Y(\i_lm[5] ));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_12 (.A(
        \write_addr[12]_net_1 ), .B(\read_addr[12]_net_1 ), .C(
        GND_net_1), .D(GND_net_1), .FCI(fifo_level_cry_11_net_1), .S(
        \fifo_level[12] ), .Y(), .FCO(fifo_level_cry_12_net_1));
    SLE \d0[21]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[21]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[17]  (.A(\state[0]_net_1 ), .B(
        \c1[17]_net_1 ), .Y(\n_HWDATA[17]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[10]  (.A(\state[0]_net_1 ), .B(
        \c1[10]_net_1 ), .Y(\n_HWDATA[10]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_RNO_1 (.A(\fifo_level[3] ), .B(
        \fifo_level[4] ), .C(\fifo_level[10] ), .D(\fifo_level[12] ), 
        .Y(m13_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(\i_cry[5]_net_1 ));
    SLE \c0[20]  (.D(din[20]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[20]_net_1 ));
    SLE \read_addr[0]  (.D(read_addr_inc_s_1_419_Y), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[0]_net_1 ));
    CFG3 #( .INIT(8'h01) )  n_d04_i_4_N_4L5 (.A(\i[4]_net_1 ), .B(
        \i[3]_net_1 ), .C(\i[5]_net_1 ), .Y(n_d04_i_4_N_4L5_net_1));
    SLE \j[1]  (.D(N_3470_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\j[1]_net_1 ));
    SLE full_ret_1 (.D(\fifo_level[12] ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\fifo_level_reto[12] ));
    ARI1 #( .INIT(20'h4AA00) )  read_addr_inc_s_13 (.A(VCC_net_1), .B(
        \read_addroi[13] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        read_addr_inc_cry_12_net_1), .S(\read_addr_inc_reti[13] ), .Y()
        , .FCO());
    CFG2 #( .INIT(4'h2) )  \state_RNIKSEJ[4]  (.A(read_en), .B(
        \state[4]_net_1 ), .Y(N_3888));
    SLE \HWDATA[22]  (.D(\n_HWDATA[22]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[22]));
    SLE \write_block_addr[13]  (.D(\next_write_addr[13] ), .CLK(mclk_1)
        , .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[13]_net_1 ));
    SLE \write_block_addr[8]  (.D(\next_write_addr[8] ), .CLK(mclk_1), 
        .EN(n_write_block_addr_0_sqmuxa), .ALn(N_4047_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\write_block_addr[8]_net_1 ));
    SLE \write_addr[7]  (.D(\next_write_addr[7] ), .CLK(mclk_1), .EN(
        N_126), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\write_addr[7]_net_1 ));
    SLE read_addr_ret_3 (.D(\read_addr_inc_reti[10] ), .CLK(mclk_1), 
        .EN(N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[10] ));
    CFG4 #( .INIT(16'h5503) )  \i_lm_0[0]  (.A(\i[0]_net_1 ), .B(
        N_3891), .C(un1_n_HWRITE_0_sqmuxa_7_0_2_net_1), .D(
        n_d04_i_RNIVD122_net_1), .Y(\i_lm[0] ));
    SLE \d0[6]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6]), .CLK(
        mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[6]));
    SLE \read_addr[9]  (.D(\read_addroi[9] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[9]_net_1 ));
    SLE \c0[28]  (.D(din[28]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[28]_net_1 ));
    SLE \addr[6]  (.D(\n_addr[6] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[6]_net_1 ));
    SLE \i[3]  (.D(\i_lm[3] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[3]_net_1 ));
    SLE \HWDATA[30]  (.D(\n_HWDATA[30]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[30]));
    CFG4 #( .INIT(16'hAA03) )  \i_lm_0[4]  (.A(\i_s[4] ), .B(N_3891), 
        .C(un1_n_HWRITE_0_sqmuxa_7_0_2_net_1), .D(
        n_d04_i_RNIVD122_net_1), .Y(\i_lm[4] ));
    CFG2 #( .INIT(4'h2) )  \HADDR_2[4]  (.A(\addr[2]_net_1 ), .B(
        test_0_HADDR[16]), .Y(test_0_HADDR[4]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[8]  (.A(\state[0]_net_1 ), .B(
        \c1[8]_net_1 ), .Y(\n_HWDATA[8]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[18]  (.A(\state[0]_net_1 ), .B(
        \c1[18]_net_1 ), .Y(\n_HWDATA[18]_net_1 ));
    SLE \HWDATA[6]  (.D(\n_HWDATA[6]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[6]));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_11 (.A(
        \write_addr[11]_net_1 ), .B(\read_addr[11]_net_1 ), .C(
        GND_net_1), .D(GND_net_1), .FCI(fifo_level_cry_10_net_1), .S(
        full_2lto11), .Y(), .FCO(fifo_level_cry_11_net_1));
    SLE \c1[16]  (.D(\c0[16]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[16]_net_1 ));
    SLE read_addr_ret (.D(\read_addr_inc_reti[13] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addroi[13] ));
    SLE \read_addr[2]  (.D(\read_addroi[2] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[2]_net_1 ));
    SLE \a_empty[0]  (.D(empty_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\a_empty[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \state_ns_x2[1]  (.A(\sync_wen[1]_net_1 ), 
        .B(\sync_wen[2]_net_1 ), .Y(N_246_i));
    CFG2 #( .INIT(4'h8) )  un1_n_HWRITE_0_sqmuxa_4_0_0_a3 (.A(
        \state[2]_net_1 ), .B(u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0)
        , .Y(N_126));
    SLE \c0[3]  (.D(din[3]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_3 (.A(VCC_net_1), 
        .B(\write_addr[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_2_net_1), .S(\next_write_addr[3] ), .Y(), 
        .FCO(next_write_addr_cry_3_net_1));
    SLE \j[0]  (.D(N_3471_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\j[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[31]  (.A(\state[0]_net_1 ), .B(
        \c1[31]_net_1 ), .Y(\n_HWDATA[31]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_9 (.A(
        \write_addr[9]_net_1 ), .B(\read_addr[9]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_8_net_1), .S(
        \fifo_level[9] ), .Y(), .FCO(fifo_level_cry_9_net_1));
    SLE \read_addr[4]  (.D(\read_addroi[4] ), .CLK(mclk_1), .EN(
        N_3845_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\read_addr[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  pipeline_cmd_RNIP2OC (.A(test_0_HADDR[16]), 
        .Y(test_0_HADDR_i_0));
    CFG3 #( .INIT(8'h80) )  n_d04_i_a3_2 (.A(\i[4]_net_1 ), .B(
        \i[3]_net_1 ), .C(\i[5]_net_1 ), .Y(N_3489));
    SLE \c1[7]  (.D(\c0[7]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c1[7]_net_1 ));
    SLE \addr[3]  (.D(\n_addr[3] ), .CLK(mclk_1), .EN(N_272_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\addr[3]_net_1 ));
    SLE \i[1]  (.D(\i_lm[1] ), .CLK(mclk_1), .EN(ie), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\i[1]_net_1 ));
    SLE \c0[16]  (.D(din[16]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[16]_net_1 ));
    SLE \HWDATA[20]  (.D(\n_HWDATA[20]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[20]));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[12]  (.A(\state[0]_net_1 ), .B(
        \c1[12]_net_1 ), .Y(\n_HWDATA[12]_net_1 ));
    SLE \HWDATA[29]  (.D(\n_HWDATA[29]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[29]));
    CFG4 #( .INIT(16'h0001) )  empty_RNO_0 (.A(\fifo_level[6] ), .B(
        \fifo_level[7] ), .C(\fifo_level[8] ), .D(\fifo_level[9] ), .Y(
        m13_5));
    CFG3 #( .INIT(8'h80) )  n_write_block_addr_0_sqmuxa_0_a3 (.A(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .B(\isl[1]_net_1 ), 
        .C(\state[2]_net_1 ), .Y(n_write_block_addr_0_sqmuxa));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[26]  (.A(\state[0]_net_1 ), .B(
        \c1[26]_net_1 ), .Y(\n_HWDATA[26]_net_1 ));
    CFG4 #( .INIT(16'h1DDD) )  full_ret_RNO_0 (.A(full_2lto11), .B(
        fifo_level_cry_10_RNIIKKL1_net_1), .C(\fifo_level[3] ), .D(
        \fifo_level[4] ), .Y(m20_1));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[11]  (.A(\state[0]_net_1 ), .B(
        \c1[11]_net_1 ), .Y(\n_HWDATA[11]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_10 (.A(
        \write_addr[10]_net_1 ), .B(\read_addr[10]_net_1 ), .C(
        GND_net_1), .D(GND_net_1), .FCI(fifo_level_cry_9_net_1), .S(
        \fifo_level[10] ), .Y(), .FCO(fifo_level_cry_10_net_1));
    SLE \a_empty[2]  (.D(\a_empty[1]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\a_empty[2]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[7]  (.A(
        \write_addr[7]_net_1 ), .B(\read_addr[7]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[7] ));
    SLE \a_full[0]  (.D(full), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\a_full[0]_net_1 ));
    SLE \c1[11]  (.D(\c0[11]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[11]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  next_write_addr_cry_6 (.A(VCC_net_1), 
        .B(\write_addr[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        next_write_addr_cry_5_net_1), .S(\next_write_addr[6] ), .Y(), 
        .FCO(next_write_addr_cry_6_net_1));
    SLE \HWDATA[9]  (.D(\n_HWDATA[9]_net_1 ), .CLK(mclk_1), .EN(
        un25_0_0_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        test_0_HWDATA[9]));
    ARI1 #( .INIT(20'h5AA55) )  fifo_level_cry_1 (.A(
        \write_addr[1]_net_1 ), .B(\read_addr[1]_net_1 ), .C(GND_net_1)
        , .D(GND_net_1), .FCI(fifo_level_cry_0_net_1), .S(
        \fifo_level[1] ), .Y(), .FCO(fifo_level_cry_1_net_1));
    SLE \c1[27]  (.D(\c0[27]_net_1 ), .CLK(mclk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\c1[27]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \n_addr_iv_0[4]  (.A(
        \write_addr[4]_net_1 ), .B(\read_addr[4]_net_1 ), .C(N_3849), 
        .D(\state[2]_net_1 ), .Y(\n_addr[4] ));
    CFG4 #( .INIT(16'hFFD5) )  n_d04_i_4 (.A(n_d04_i_4_N_3L3_net_1), 
        .B(n_d04_i_4_N_4L5_net_1), .C(N_3474), .D(
        n_d04_i_4_N_2L1_net_1), .Y(n_d04_i_4_net_1));
    CFG3 #( .INIT(8'hFE) )  n_d04_i (.A(N_3484), .B(n_d04_i_4_net_1), 
        .C(N_3489), .Y(N_3467));
    SLE \d0[30]  (.D(u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30]), 
        .CLK(mclk_1), .EN(N_3847_i), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dout[30]));
    CFG4 #( .INIT(16'hFFF8) )  n_d04_i_a3_RNISQ4N6 (.A(
        un1_n_HWRITE_1_sqmuxa_2_i_0_233_i_o3_i_o2_d), .B(
        un1_n_HWRITE_1_sqmuxa_2_i_0_i_o3_i_o2_0_4), .C(ilde_0_1), .D(
        N_3886), .Y(ie));
    SLE full_ret (.D(N_36_mux), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(N_36_mux_reto));
    CFG2 #( .INIT(4'h4) )  \n_HWDATA[25]  (.A(\state[0]_net_1 ), .B(
        \c1[25]_net_1 ), .Y(\n_HWDATA[25]_net_1 ));
    SLE \c0[11]  (.D(din[11]), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\c0[11]_net_1 ));
    
endmodule


module sync_logic_1s_2(
       status_0,
       almost_full_sync,
       sdclk_n_1,
       mclk_1,
       N_4047_i
    );
input  status_0;
output almost_full_sync;
input  sdclk_n_1;
input  mclk_1;
input  N_4047_i;

    wire \update_ack_dly[1]_net_1 , \update_ack_dly_i[1] , 
        \update_strobe_dly[1]_net_1 , VCC_net_1, 
        \update_strobe_dly[0]_net_1 , GND_net_1, 
        \update_strobe_dly[2]_net_1 , \update_strobe_dly[3]_net_1 , 
        update_strobe_net_1, update_ack_net_1, \data_buf[0]_net_1 , 
        un1_update_strobe_dly_1, data_buf6_i_net_1, 
        \update_ack_dly[0]_net_1 ;
    
    SLE update_strobe (.D(\update_ack_dly_i[1] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(update_strobe_net_1));
    GND GND (.Y(GND_net_1));
    SLE \data_buf_sync[0]  (.D(\data_buf[0]_net_1 ), .CLK(mclk_1), .EN(
        un1_update_strobe_dly_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        almost_full_sync));
    CFG2 #( .INIT(4'h9) )  data_buf6_i (.A(update_strobe_net_1), .B(
        \update_ack_dly[1]_net_1 ), .Y(data_buf6_i_net_1));
    SLE \data_buf[0]  (.D(status_0), .CLK(sdclk_n_1), .EN(
        data_buf6_i_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_buf[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  update_strobe_RNO (.A(
        \update_ack_dly[1]_net_1 ), .Y(\update_ack_dly_i[1] ));
    SLE \update_ack_dly[1]  (.D(\update_ack_dly[0]_net_1 ), .CLK(
        sdclk_n_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[1]_net_1 ));
    SLE \update_strobe_dly[2]  (.D(\update_strobe_dly[1]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[2]_net_1 ));
    SLE \update_strobe_dly[0]  (.D(update_strobe_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[0]_net_1 ));
    SLE \update_strobe_dly[3]  (.D(\update_strobe_dly[2]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[3]_net_1 ));
    SLE \update_ack_dly[0]  (.D(update_ack_net_1), .CLK(sdclk_n_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[0]_net_1 ));
    SLE update_ack (.D(\update_strobe_dly[3]_net_1 ), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        update_ack_net_1));
    CFG2 #( .INIT(4'h6) )  un1_update_strobe_dly (.A(update_ack_net_1), 
        .B(\update_strobe_dly[3]_net_1 ), .Y(un1_update_strobe_dly_1));
    SLE \update_strobe_dly[1]  (.D(\update_strobe_dly[0]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[1]_net_1 ));
    
endmodule


module sync_logic_1s(
       un1_ctrl,
       sdctrl_start_i2s,
       sdclk_n_1,
       mclk_1,
       N_4047_i
    );
input  un1_ctrl;
output sdctrl_start_i2s;
input  sdclk_n_1;
input  mclk_1;
input  N_4047_i;

    wire \update_ack_dly[1]_net_1 , \update_ack_dly_i[1] , 
        \update_strobe_dly[1]_net_1 , VCC_net_1, 
        \update_strobe_dly[0]_net_1 , GND_net_1, 
        \update_strobe_dly[2]_net_1 , \update_strobe_dly[3]_net_1 , 
        update_strobe_net_1, update_ack_net_1, \data_buf[0]_net_1 , 
        un1_update_strobe_dly_net_1, data_buf6_i_net_1, 
        \update_ack_dly[0]_net_1 ;
    
    SLE update_strobe (.D(\update_ack_dly_i[1] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(update_strobe_net_1));
    GND GND (.Y(GND_net_1));
    SLE \data_buf_sync[0]  (.D(\data_buf[0]_net_1 ), .CLK(mclk_1), .EN(
        un1_update_strobe_dly_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdctrl_start_i2s));
    CFG2 #( .INIT(4'h9) )  data_buf6_i (.A(update_strobe_net_1), .B(
        \update_ack_dly[1]_net_1 ), .Y(data_buf6_i_net_1));
    SLE \data_buf[0]  (.D(un1_ctrl), .CLK(sdclk_n_1), .EN(
        data_buf6_i_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_buf[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  update_strobe_RNO (.A(
        \update_ack_dly[1]_net_1 ), .Y(\update_ack_dly_i[1] ));
    SLE \update_ack_dly[1]  (.D(\update_ack_dly[0]_net_1 ), .CLK(
        sdclk_n_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[1]_net_1 ));
    SLE \update_strobe_dly[2]  (.D(\update_strobe_dly[1]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[2]_net_1 ));
    SLE \update_strobe_dly[0]  (.D(update_strobe_net_1), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[0]_net_1 ));
    SLE \update_strobe_dly[3]  (.D(\update_strobe_dly[2]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[3]_net_1 ));
    SLE \update_ack_dly[0]  (.D(update_ack_net_1), .CLK(sdclk_n_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_ack_dly[0]_net_1 ));
    SLE update_ack (.D(\update_strobe_dly[3]_net_1 ), .CLK(mclk_1), 
        .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        update_ack_net_1));
    CFG2 #( .INIT(4'h6) )  un1_update_strobe_dly (.A(update_ack_net_1), 
        .B(\update_strobe_dly[3]_net_1 ), .Y(
        un1_update_strobe_dly_net_1));
    SLE \update_strobe_dly[1]  (.D(\update_strobe_dly[0]_net_1 ), .CLK(
        mclk_1), .EN(VCC_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \update_strobe_dly[1]_net_1 ));
    
endmodule


module mem_controller(
       din,
       status,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0,
       test_0_HWDATA,
       test_0_HADDR,
       source_right,
       source_left,
       dsd138_ctrl,
       test_0_HADDR_i_0,
       test_0_HTRANS_0,
       state_0_d0,
       state_0_0,
       bus_state_0,
       sound_card_ctrl_7,
       sound_card_ctrl_6,
       sound_card_ctrl_5,
       sound_card_ctrl_0,
       sound_card_ctrl_1,
       sound_card_ctrl_2,
       cnt_0,
       is_last_data,
       test_0_HWRITE,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       wen,
       buffer_under_runlde_0_a6_2,
       sdclk_n_1,
       in_bck_1,
       master_lrck,
       use_dsd,
       i2s_start,
       mclk_1,
       N_4047_i
    );
input  [31:0] din;
output [7:6] status;
input  [31:0] u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0;
output [31:0] test_0_HWDATA;
output [16:2] test_0_HADDR;
output [31:0] source_right;
output [31:0] source_left;
output [2:0] dsd138_ctrl;
output test_0_HADDR_i_0;
output test_0_HTRANS_0;
input  state_0_d0;
input  state_0_0;
input  bus_state_0;
input  sound_card_ctrl_7;
input  sound_card_ctrl_6;
input  sound_card_ctrl_5;
input  sound_card_ctrl_0;
input  sound_card_ctrl_1;
input  sound_card_ctrl_2;
input  cnt_0;
input  is_last_data;
output test_0_HWRITE;
input  u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
input  wen;
output buffer_under_runlde_0_a6_2;
input  sdclk_n_1;
input  in_bck_1;
input  master_lrck;
output use_dsd;
output i2s_start;
input  mclk_1;
input  N_4047_i;

    wire \k[2]_net_1 , VCC_net_1, k_n2_net_1, ke, GND_net_1, 
        \k[3]_net_1 , k_n3_net_1, \k[4]_net_1 , k_n4_net_1, 
        \k[0]_net_1 , N_1270, \k[1]_net_1 , k_n1_net_1, 
        \pcm_left_RNO[28]_net_1 , un1_state_6_i, N_1257_i, 
        \pcm_left_RNO[30]_net_1 , N_1237_i, \sdctrl_bck_divider[0] , 
        N_3826_i, \sdctrl_bck_divider[1] , \sdctrl_bck_divider[2] , 
        N_1229_i, \pcm_left_RNO[14]_net_1 , N_1209_i, 
        \pcm_left_RNO[16]_net_1 , N_1189_i, \pcm_left_RNO[18]_net_1 , 
        N_1169_i, \pcm_left_RNO[20]_net_1 , N_1149_i, 
        \pcm_left_RNO[22]_net_1 , N_1129_i, \pcm_left_RNO[24]_net_1 , 
        N_1109_i, \pcm_left_RNO[26]_net_1 , N_1089_i, \left[30]_net_1 , 
        \dout[30] , un1_state_7_i_a3_2_net_1, \left[31]_net_1 , 
        \dout[31] , \pcm_left_RNO[0]_net_1 , N_1069_i, 
        \pcm_left_RNO[2]_net_1 , N_1049_i, \pcm_left_RNO[4]_net_1 , 
        N_1029_i, \pcm_left_RNO[6]_net_1 , N_1009_i, 
        \pcm_left_RNO[8]_net_1 , N_989_i, \pcm_left_RNO[10]_net_1 , 
        N_969_i, \pcm_left_RNO[12]_net_1 , \left[15]_net_1 , 
        \dout[15] , \left[16]_net_1 , \dout[16] , \left[17]_net_1 , 
        \dout[17] , \left[18]_net_1 , \dout[18] , \left[19]_net_1 , 
        \dout[19] , \left[20]_net_1 , \dout[20] , \left[21]_net_1 , 
        \dout[21] , \left[22]_net_1 , \dout[22] , \left[23]_net_1 , 
        \dout[23] , \left[24]_net_1 , \dout[24] , \left[25]_net_1 , 
        \dout[25] , \left[26]_net_1 , \dout[26] , \left[27]_net_1 , 
        \dout[27] , \left[28]_net_1 , \dout[28] , \left[29]_net_1 , 
        \dout[29] , \left[0]_net_1 , \dout[0] , \left[1]_net_1 , 
        \dout[1] , \left[2]_net_1 , \dout[2] , \left[3]_net_1 , 
        \dout[3] , \left[4]_net_1 , \dout[4] , \left[5]_net_1 , 
        \dout[5] , \left[6]_net_1 , \dout[6] , \left[7]_net_1 , 
        \dout[7] , \left[8]_net_1 , \dout[8] , \left[9]_net_1 , 
        \dout[9] , \left[10]_net_1 , \dout[10] , \left[11]_net_1 , 
        \dout[11] , \left[12]_net_1 , \dout[12] , \left[13]_net_1 , 
        \dout[13] , \left[14]_net_1 , \dout[14] , N_949_i, 
        \pcm_right_RNO[18]_net_1 , N_929_i, \pcm_right_RNO[20]_net_1 , 
        N_909_i, \pcm_right_RNO[22]_net_1 , N_889_i, 
        \pcm_right_RNO[24]_net_1 , N_869_i, \pcm_right_RNO[26]_net_1 , 
        N_849_i, \pcm_right_RNO[28]_net_1 , N_829_i, 
        \pcm_right_RNO[30]_net_1 , N_809_i, \pcm_right_RNO[2]_net_1 , 
        N_789_i, \pcm_right_RNO[4]_net_1 , N_769_i, 
        \pcm_right_RNO[6]_net_1 , N_749_i, \pcm_right_RNO[8]_net_1 , 
        N_729_i, \pcm_right_RNO[10]_net_1 , N_709_i, 
        \pcm_right_RNO[12]_net_1 , N_689_i, N_679, N_669_i, N_659, 
        \pcm_right_RNO[0]_net_1 , N_637_i, flag_net_1, flag_ldmx_net_1, 
        N_3842_i, N_3820_i, N_3822_i, sdctrl_use_dsd, read_en_net_1, 
        N_9_i, \state[0]_net_1 , N_9_i_0, \state[1]_net_1 , m10_i, 
        old_lrck_net_1, old_bck_net_1, N_166, N_3843, n_pcm13_0_net_1, 
        k_n0_0_875_a3_0_0_net_1, N_3825, N_175, N_3829, un1_ctrl_net_1, 
        N_162, un1_state_7_i_a3_1_net_1, k_c2_net_1, sdctrl_start_i2s, 
        almost_full_sync, \pcm_dec[1] , N_3833, m8_0_0, m8_0_0_0, 
        flag_en_net_1, m8_0_2;
    
    CFG4 #( .INIT(16'h8000) )  n_pcm13 (.A(\k[0]_net_1 ), .B(
        n_pcm13_0_net_1), .C(\k[2]_net_1 ), .D(\k[1]_net_1 ), .Y(N_175)
        );
    SLE \pcm_left[22]  (.D(\pcm_left_RNO[22]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[22]));
    SLE \state[0]  (.D(N_9_i_0), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[25]  (.A(\state[1]_net_1 ), 
        .B(\dout[25] ), .Y(N_869_i));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[17]  (.A(\state[1]_net_1 ), 
        .B(\left[17]_net_1 ), .Y(N_1189_i));
    SLE \pcm_right[9]  (.D(N_729_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[9]));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[29]  (.A(\state[1]_net_1 ), 
        .B(\left[29]_net_1 ), .Y(N_1257_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[2]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[2]_net_1 ), .Y(\pcm_left_RNO[2]_net_1 ));
    SLE \left[9]  (.D(\dout[9] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[9]_net_1 ));
    SLE \pcm_left[27]  (.D(N_1089_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[27]));
    CFG4 #( .INIT(16'h48C0) )  k_n2 (.A(\k[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(\k[2]_net_1 ), .D(\k[1]_net_1 ), .Y(
        k_n2_net_1));
    CFG4 #( .INIT(16'h3307) )  \n_read_en.m8_0_0  (.A(almost_full_sync)
        , .B(sdctrl_start_i2s), .C(\state[0]_net_1 ), .D(
        \state[1]_net_1 ), .Y(m8_0_0));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[23]  (.A(\state[1]_net_1 ), 
        .B(\dout[23] ), .Y(N_889_i));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[5]  (.A(\state[1]_net_1 ), .B(
        \left[5]_net_1 ), .Y(N_1029_i));
    SLE \pcm_right[20]  (.D(\pcm_right_RNO[20]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[20]));
    SLE \pcm_left[9]  (.D(N_989_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[9]));
    SLE \k[1]  (.D(k_n1_net_1), .CLK(mclk_1), .EN(ke), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\k[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[10]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[10] ), .Y(\pcm_right_RNO[10]_net_1 ));
    SLE \pcm_left[14]  (.D(\pcm_left_RNO[14]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[14]));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[16]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[16] ), .Y(N_659));
    SLE \pcm_right[24]  (.D(\pcm_right_RNO[24]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[24]));
    SLE \pcm_left[26]  (.D(\pcm_left_RNO[26]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[26]));
    SLE \pcm_right[11]  (.D(N_709_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[11]));
    SLE \bck_divider[2]  (.D(\sdctrl_bck_divider[2] ), .CLK(mclk_1), 
        .EN(N_3826_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(dsd138_ctrl[2]));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[14]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[14] ), .Y(N_679));
    CFG2 #( .INIT(4'h8) )  n_pcm13_0 (.A(\k[3]_net_1 ), .B(
        \k[4]_net_1 ), .Y(n_pcm13_0_net_1));
    SLE \pcm_right[0]  (.D(\pcm_right_RNO[0]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[0]));
    SLE flag (.D(flag_ldmx_net_1), .CLK(mclk_1), .EN(N_3842_i), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(flag_net_1));
    CFG4 #( .INIT(16'h4000) )  pcm_dec_1 (.A(\k[0]_net_1 ), .B(
        n_pcm13_0_net_1), .C(\k[2]_net_1 ), .D(\k[1]_net_1 ), .Y(
        \pcm_dec[1] ));
    CFG4 #( .INIT(16'h60A0) )  k_n4 (.A(\k[4]_net_1 ), .B(\k[3]_net_1 )
        , .C(\state[1]_net_1 ), .D(k_c2_net_1), .Y(k_n4_net_1));
    SLE \left[6]  (.D(\dout[6] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[6]_net_1 ));
    SLE \left[20]  (.D(\dout[20] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[20]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[5]  (.A(\state[1]_net_1 ), 
        .B(\dout[5] ), .Y(N_769_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[12]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[12] ), .Y(\pcm_right_RNO[12]_net_1 ));
    CFG4 #( .INIT(16'hE6A2) )  n_k10_RNIAL0F1 (.A(\state[1]_net_1 ), 
        .B(\state[0]_net_1 ), .C(N_162), .D(N_166), .Y(ke));
    SLE \pcm_right[25]  (.D(N_869_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[25]));
    sync_logic_1s_1 usync101 (.sound_card_ctrl_0(sound_card_ctrl_5), 
        .sdctrl_use_dsd(sdctrl_use_dsd), .sdclk_n_1(sdclk_n_1), 
        .mclk_1(mclk_1), .N_4047_i(N_4047_i));
    SLE \left[19]  (.D(\dout[19] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[19]_net_1 ));
    SLE \left[12]  (.D(\dout[12] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[12]_net_1 ));
    SLE \pcm_right[1]  (.D(N_637_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[1]));
    SLE \pcm_right[31]  (.D(N_809_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[31]));
    SLE \pcm_left[6]  (.D(\pcm_left_RNO[6]_net_1 ), .CLK(mclk_1), .EN(
        un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(source_left[6])
        );
    SLE \left[18]  (.D(\dout[18] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[18]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \pcm_right[5]  (.D(N_769_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[5]));
    CFG4 #( .INIT(16'h3F07) )  \state_ns_1_0_.m8_0_0  (.A(
        almost_full_sync), .B(sdctrl_start_i2s), .C(\state[0]_net_1 ), 
        .D(\state[1]_net_1 ), .Y(m8_0_0_0));
    SLE read_en (.D(N_9_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(read_en_net_1));
    CFG4 #( .INIT(16'hFD31) )  flag_en (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(N_166), .D(N_175), .Y(flag_en_net_1));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[20]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[20] ), .Y(\pcm_right_RNO[20]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[26]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[26] ), .Y(\pcm_right_RNO[26]_net_1 ));
    SLE use_dsd_inst_1 (.D(sdctrl_use_dsd), .CLK(mclk_1), .EN(N_3826_i)
        , .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(use_dsd));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[12]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[12]_net_1 ), .Y(\pcm_left_RNO[12]_net_1 )
        );
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[7]  (.A(\state[1]_net_1 ), 
        .B(\dout[7] ), .Y(N_749_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[24]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[24] ), .Y(\pcm_right_RNO[24]_net_1 ));
    SLE \pcm_left[24]  (.D(\pcm_left_RNO[24]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[24]));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[1]  (.A(\state[1]_net_1 ), .B(
        \left[1]_net_1 ), .Y(N_1069_i));
    CFG2 #( .INIT(4'h8) )  un1_ctrl (.A(sound_card_ctrl_7), .B(
        sound_card_ctrl_6), .Y(un1_ctrl_net_1));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[24]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[24]_net_1 ), .Y(\pcm_left_RNO[24]_net_1 )
        );
    SLE \left[4]  (.D(\dout[4] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[4]_net_1 ));
    SLE \left[16]  (.D(\dout[16] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[16]_net_1 ));
    SLE \k[4]  (.D(k_n4_net_1), .CLK(mclk_1), .EN(ke), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\k[4]_net_1 ));
    SLE \pcm_right[28]  (.D(\pcm_right_RNO[28]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[28]));
    SLE \left[2]  (.D(\dout[2] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[2]_net_1 ));
    SLE \pcm_right[29]  (.D(N_829_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[29]));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[22]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[22] ), .Y(\pcm_right_RNO[22]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[20]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[20]_net_1 ), .Y(\pcm_left_RNO[20]_net_1 )
        );
    CFG3 #( .INIT(8'h20) )  n_k10_RNI7O731 (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(N_166), .Y(N_3843));
    SLE \left[29]  (.D(\dout[29] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[29]_net_1 ));
    SLE \left[22]  (.D(\dout[22] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[22]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[6]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[6]_net_1 ), .Y(\pcm_left_RNO[6]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[26]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[26]_net_1 ), .Y(\pcm_left_RNO[26]_net_1 )
        );
    SLE \pcm_right[16]  (.D(N_659), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[16]));
    SLE \k[2]  (.D(k_n2_net_1), .CLK(mclk_1), .EN(ke), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\k[2]_net_1 ));
    SLE \pcm_right[6]  (.D(\pcm_right_RNO[6]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[6]));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[13]  (.A(\state[1]_net_1 ), 
        .B(\left[13]_net_1 ), .Y(N_1229_i));
    SLE \left[28]  (.D(\dout[28] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[28]_net_1 ));
    SLE \pcm_left[2]  (.D(\pcm_left_RNO[2]_net_1 ), .CLK(mclk_1), .EN(
        un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(source_left[2])
        );
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[21]  (.A(\state[1]_net_1 ), 
        .B(\left[21]_net_1 ), .Y(N_1149_i));
    VCC VCC (.Y(VCC_net_1));
    sync_logic_3s usync102 (.sound_card_ctrl({sound_card_ctrl_2, 
        sound_card_ctrl_1, sound_card_ctrl_0}), .sdctrl_bck_divider({
        \sdctrl_bck_divider[2] , \sdctrl_bck_divider[1] , 
        \sdctrl_bck_divider[0] }), .mclk_1(mclk_1), .sdclk_n_1(
        sdclk_n_1), .N_4047_i(N_4047_i));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[9]  (.A(\state[1]_net_1 ), 
        .B(\dout[9] ), .Y(N_729_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[18]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[18] ), .Y(\pcm_right_RNO[18]_net_1 ));
    SLE \pcm_left[7]  (.D(N_1009_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[7]));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[15]  (.A(\state[1]_net_1 ), 
        .B(\left[15]_net_1 ), .Y(N_1209_i));
    SLE \pcm_right[27]  (.D(N_849_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[27]));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[18]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[18]_net_1 ), .Y(\pcm_left_RNO[18]_net_1 )
        );
    SLE \left[26]  (.D(\dout[26] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[26]_net_1 ));
    SLE \pcm_right[8]  (.D(\pcm_right_RNO[8]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[8]));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[30]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[30] ), .Y(\pcm_right_RNO[30]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[6]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[6] ), .Y(\pcm_right_RNO[6]_net_1 ));
    SLE \pcm_left[10]  (.D(\pcm_left_RNO[10]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[10]));
    CFG3 #( .INIT(8'h80) )  k_c2 (.A(\k[2]_net_1 ), .B(\k[1]_net_1 ), 
        .C(\k[0]_net_1 ), .Y(k_c2_net_1));
    CFG3 #( .INIT(8'h53) )  sound_card_start_RNO (.A(sdctrl_start_i2s), 
        .B(\state[0]_net_1 ), .C(\state[1]_net_1 ), .Y(N_3822_i));
    SLE \pcm_right[23]  (.D(N_889_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[23]));
    CFG4 #( .INIT(16'h1D15) )  un1_state_6_0_o2_1_RNIPOT91 (.A(
        \state[0]_net_1 ), .B(\state[1]_net_1 ), .C(N_3829), .D(N_162), 
        .Y(un1_state_6_i));
    CFG2 #( .INIT(4'h7) )  un1_state_6_0_o2_1 (.A(N_175), .B(
        flag_net_1), .Y(N_3829));
    SLE \pcm_right[22]  (.D(\pcm_right_RNO[22]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[22]));
    CFG2 #( .INIT(4'h8) )  \n_read_en.N_3820_i  (.A(sdctrl_start_i2s), 
        .B(almost_full_sync), .Y(N_3820_i));
    SLE \k[3]  (.D(k_n3_net_1), .CLK(mclk_1), .EN(ke), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\k[3]_net_1 ));
    SLE \k[0]  (.D(N_1270), .CLK(mclk_1), .EN(ke), .ALn(N_4047_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\k[0]_net_1 ));
    SLE \bck_divider[1]  (.D(\sdctrl_bck_divider[1] ), .CLK(mclk_1), 
        .EN(N_3826_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(dsd138_ctrl[1]));
    SLE \pcm_left[30]  (.D(\pcm_left_RNO[30]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[30]));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[4]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[4] ), .Y(\pcm_right_RNO[4]_net_1 ));
    SLE \left[5]  (.D(\dout[5] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[5]_net_1 ));
    SLE \left[1]  (.D(\dout[1] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[1]_net_1 ));
    SLE \left[14]  (.D(\dout[14] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[14]_net_1 ));
    SLE \pcm_right[2]  (.D(\pcm_right_RNO[2]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[2]));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[19]  (.A(\state[1]_net_1 ), 
        .B(\left[19]_net_1 ), .Y(N_1169_i));
    SLE \pcm_left[0]  (.D(\pcm_left_RNO[0]_net_1 ), .CLK(mclk_1), .EN(
        un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(source_left[0])
        );
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[28]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[28] ), .Y(\pcm_right_RNO[28]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[11]  (.A(\state[1]_net_1 ), 
        .B(\dout[11] ), .Y(N_709_i));
    CFG2 #( .INIT(4'hB) )  un1_state_6_0_o2_0 (.A(\state[1]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(N_3825));
    SLE \left[8]  (.D(\dout[8] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[8]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[27]  (.A(\state[1]_net_1 ), 
        .B(\left[27]_net_1 ), .Y(N_1089_i));
    SLE \pcm_left[19]  (.D(N_1169_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[19]));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[17]  (.A(\state[1]_net_1 ), 
        .B(\dout[17] ), .Y(N_949_i));
    SLE \left[7]  (.D(\dout[7] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[7]_net_1 ));
    CFG3 #( .INIT(8'h08) )  un1_state_7_i_a3_1 (.A(\state[1]_net_1 ), 
        .B(N_175), .C(flag_net_1), .Y(un1_state_7_i_a3_1_net_1));
    SLE \pcm_right[21]  (.D(N_909_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[21]));
    SLE \pcm_right[10]  (.D(\pcm_right_RNO[10]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[10]));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[0]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[0]_net_1 ), .Y(\pcm_left_RNO[0]_net_1 ));
    SLE \left[31]  (.D(\dout[31] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[31]_net_1 ));
    SLE \left[0]  (.D(\dout[0] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[0]_net_1 ));
    SLE \pcm_right[14]  (.D(N_679), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[14]));
    SLE \pcm_left[20]  (.D(\pcm_left_RNO[20]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[20]));
    SLE \pcm_left[18]  (.D(\pcm_left_RNO[18]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[18]));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[1]  (.A(\state[1]_net_1 ), 
        .B(\dout[1] ), .Y(N_637_i));
    SLE \left[17]  (.D(\dout[17] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[17]_net_1 ));
    SLE \left[24]  (.D(\dout[24] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[24]_net_1 ));
    SLE \bck_divider[0]  (.D(\sdctrl_bck_divider[0] ), .CLK(mclk_1), 
        .EN(N_3826_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(dsd138_ctrl[0]));
    CFG3 #( .INIT(8'hEC) )  \state_ns_1_0_.m10_i  (.A(\state[1]_net_1 )
        , .B(N_3843), .C(sdctrl_start_i2s), .Y(m10_i));
    SLE \pcm_left[15]  (.D(N_1209_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[15]));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[8]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[8]_net_1 ), .Y(\pcm_left_RNO[8]_net_1 ));
    SLE \left[15]  (.D(\dout[15] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[15]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[19]  (.A(\state[1]_net_1 ), 
        .B(\dout[19] ), .Y(N_929_i));
    SLE \pcm_right[15]  (.D(N_669_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[15]));
    CFG4 #( .INIT(16'h00F7) )  \n_read_en.N_9_i  (.A(\state[0]_net_1 ), 
        .B(\state[1]_net_1 ), .C(N_162), .D(m8_0_2), .Y(N_9_i));
    bigfifo ufifo (.test_0_HADDR({test_0_HADDR[16], test_0_HADDR[15], 
        test_0_HADDR[14], test_0_HADDR[13], test_0_HADDR[12], 
        test_0_HADDR[11], test_0_HADDR[10], test_0_HADDR[9], 
        test_0_HADDR[8], test_0_HADDR[7], test_0_HADDR[6], 
        test_0_HADDR[5], test_0_HADDR[4], test_0_HADDR[3], 
        test_0_HADDR[2]}), .test_0_HWDATA({test_0_HWDATA[31], 
        test_0_HWDATA[30], test_0_HWDATA[29], test_0_HWDATA[28], 
        test_0_HWDATA[27], test_0_HWDATA[26], test_0_HWDATA[25], 
        test_0_HWDATA[24], test_0_HWDATA[23], test_0_HWDATA[22], 
        test_0_HWDATA[21], test_0_HWDATA[20], test_0_HWDATA[19], 
        test_0_HWDATA[18], test_0_HWDATA[17], test_0_HWDATA[16], 
        test_0_HWDATA[15], test_0_HWDATA[14], test_0_HWDATA[13], 
        test_0_HWDATA[12], test_0_HWDATA[11], test_0_HWDATA[10], 
        test_0_HWDATA[9], test_0_HWDATA[8], test_0_HWDATA[7], 
        test_0_HWDATA[6], test_0_HWDATA[5], test_0_HWDATA[4], 
        test_0_HWDATA[3], test_0_HWDATA[2], test_0_HWDATA[1], 
        test_0_HWDATA[0]}), .u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0({
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0]}), .dout({
        \dout[31] , \dout[30] , \dout[29] , \dout[28] , \dout[27] , 
        \dout[26] , \dout[25] , \dout[24] , \dout[23] , \dout[22] , 
        \dout[21] , \dout[20] , \dout[19] , \dout[18] , \dout[17] , 
        \dout[16] , \dout[15] , \dout[14] , \dout[13] , \dout[12] , 
        \dout[11] , \dout[10] , \dout[9] , \dout[8] , \dout[7] , 
        \dout[6] , \dout[5] , \dout[4] , \dout[3] , \dout[2] , 
        \dout[1] , \dout[0] }), .status({status[7], status[6]}), .din({
        din[31], din[30], din[29], din[28], din[27], din[26], din[25], 
        din[24], din[23], din[22], din[21], din[20], din[19], din[18], 
        din[17], din[16], din[15], din[14], din[13], din[12], din[11], 
        din[10], din[9], din[8], din[7], din[6], din[5], din[4], 
        din[3], din[2], din[1], din[0]}), .bus_state_0(bus_state_0), 
        .state_0_0(state_0_0), .state_0_d0(state_0_d0), 
        .test_0_HTRANS_0(test_0_HTRANS_0), .test_0_HADDR_i_0(
        test_0_HADDR_i_0), .buffer_under_runlde_0_a6_2(
        buffer_under_runlde_0_a6_2), .wen(wen), .read_en(read_en_net_1)
        , .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .test_0_HWRITE(
        test_0_HWRITE), .sdclk_n_1(sdclk_n_1), .is_last_data(
        is_last_data), .N_4047_i(N_4047_i), .mclk_1(mclk_1));
    SLE \pcm_left[1]  (.D(N_1069_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[1]));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[21]  (.A(\state[1]_net_1 ), 
        .B(\dout[21] ), .Y(N_909_i));
    SLE \pcm_right[30]  (.D(\pcm_right_RNO[30]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[30]));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[4]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[4]_net_1 ), .Y(\pcm_left_RNO[4]_net_1 ));
    CFG4 #( .INIT(16'h1555) )  \state_ns_1_0_.N_9_i  (.A(m8_0_0_0), .B(
        N_3843), .C(\sdctrl_bck_divider[0] ), .D(
        k_n0_0_875_a3_0_0_net_1), .Y(N_9_i_0));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[27]  (.A(\state[1]_net_1 ), 
        .B(\dout[27] ), .Y(N_849_i));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[3]  (.A(\state[1]_net_1 ), .B(
        \left[3]_net_1 ), .Y(N_1049_i));
    SLE \pcm_left[29]  (.D(N_1257_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[29]));
    SLE old_lrck (.D(master_lrck), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(old_lrck_net_1));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[0]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[0] ), .Y(\pcm_right_RNO[0]_net_1 ));
    CFG4 #( .INIT(16'hFCDC) )  un1_state_7_i_a3_2 (.A(\state[0]_net_1 )
        , .B(N_3843), .C(un1_state_7_i_a3_1_net_1), .D(N_162), .Y(
        un1_state_7_i_a3_2_net_1));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[30]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[30]_net_1 ), .Y(\pcm_left_RNO[30]_net_1 )
        );
    CFG2 #( .INIT(4'h1) )  \state_RNI5SEN[0]  (.A(\state[1]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(N_3826_i));
    SLE \left[13]  (.D(\dout[13] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[13]_net_1 ));
    SLE \pcm_left[8]  (.D(\pcm_left_RNO[8]_net_1 ), .CLK(mclk_1), .EN(
        un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(source_left[8])
        );
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[3]  (.A(\state[1]_net_1 ), 
        .B(\dout[3] ), .Y(N_789_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[14]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[14]_net_1 ), .Y(\pcm_left_RNO[14]_net_1 )
        );
    sync_logic_1s_2 usync600 (.status_0(status[7]), .almost_full_sync(
        almost_full_sync), .sdclk_n_1(sdclk_n_1), .mclk_1(mclk_1), 
        .N_4047_i(N_4047_i));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[7]  (.A(\state[1]_net_1 ), .B(
        \left[7]_net_1 ), .Y(N_1009_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[22]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[22]_net_1 ), .Y(\pcm_left_RNO[22]_net_1 )
        );
    CFG4 #( .INIT(16'hFFF1) )  \n_read_en.m8_0_2  (.A(N_166), .B(
        N_3825), .C(m8_0_0), .D(N_3833), .Y(m8_0_2));
    SLE \left[27]  (.D(\dout[27] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[27]_net_1 ));
    SLE \left[11]  (.D(\dout[11] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[11]_net_1 ));
    SLE \pcm_left[11]  (.D(N_969_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[11]));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[10]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[10]_net_1 ), .Y(\pcm_left_RNO[10]_net_1 )
        );
    SLE \pcm_left[28]  (.D(\pcm_left_RNO[28]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[28]));
    SLE \state[1]  (.D(m10_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    SLE \left[25]  (.D(\dout[25] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[25]_net_1 ));
    CFG4 #( .INIT(16'h028A) )  \n_read_en.m8_0_a3  (.A(
        \state[1]_net_1 ), .B(\state[0]_net_1 ), .C(N_175), .D(
        \pcm_dec[1] ), .Y(N_3833));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[31]  (.A(\state[1]_net_1 ), 
        .B(\left[31]_net_1 ), .Y(N_1237_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[16]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[16]_net_1 ), .Y(\pcm_left_RNO[16]_net_1 )
        );
    SLE \pcm_right[26]  (.D(\pcm_right_RNO[26]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[26]));
    SLE \pcm_right[18]  (.D(\pcm_right_RNO[18]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[18]));
    SLE \pcm_right[19]  (.D(N_929_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[19]));
    SLE \pcm_left[31]  (.D(N_1237_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[31]));
    SLE \pcm_left[5]  (.D(N_1029_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[5]));
    SLE \pcm_left[25]  (.D(N_1109_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[25]));
    SLE \pcm_left[13]  (.D(N_1229_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[13]));
    SLE \left[30]  (.D(\dout[30] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[30]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[29]  (.A(\state[1]_net_1 ), 
        .B(\dout[29] ), .Y(N_829_i));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[11]  (.A(\state[1]_net_1 ), 
        .B(\left[11]_net_1 ), .Y(N_969_i));
    SLE \pcm_left[12]  (.D(\pcm_left_RNO[12]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[12]));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[23]  (.A(\state[1]_net_1 ), 
        .B(\left[23]_net_1 ), .Y(N_1129_i));
    CFG4 #( .INIT(16'h33A0) )  k_n0_0_875 (.A(\sdctrl_bck_divider[0] ), 
        .B(\k[0]_net_1 ), .C(k_n0_0_875_a3_0_0_net_1), .D(
        \state[1]_net_1 ), .Y(N_1270));
    SLE \pcm_left[3]  (.D(N_1049_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[3]));
    SLE \pcm_right[3]  (.D(N_789_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[3]));
    SLE \left[23]  (.D(\dout[23] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[23]_net_1 ));
    CFG2 #( .INIT(4'h4) )  k_n0_0_875_a3_0_0 (.A(
        \sdctrl_bck_divider[1] ), .B(\sdctrl_bck_divider[2] ), .Y(
        k_n0_0_875_a3_0_0_net_1));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[15]  (.A(\state[1]_net_1 ), 
        .B(\dout[15] ), .Y(N_669_i));
    SLE \pcm_left[17]  (.D(N_1189_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[17]));
    CFG3 #( .INIT(8'h8A) )  n_k10 (.A(old_lrck_net_1), .B(cnt_0), .C(
        i2s_start), .Y(N_166));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[8]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[8] ), .Y(\pcm_right_RNO[8]_net_1 ));
    SLE old_bck (.D(in_bck_1), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(old_bck_net_1));
    CFG3 #( .INIT(8'hDF) )  flag_RNO (.A(\state[1]_net_1 ), .B(N_162), 
        .C(\state[0]_net_1 ), .Y(N_3842_i));
    CFG3 #( .INIT(8'hE4) )  \pcm_right_RNO[2]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\dout[2] ), .Y(\pcm_right_RNO[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[25]  (.A(\state[1]_net_1 ), 
        .B(\left[25]_net_1 ), .Y(N_1109_i));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[31]  (.A(\state[1]_net_1 ), 
        .B(\dout[31] ), .Y(N_809_i));
    CFG2 #( .INIT(4'h8) )  \pcm_right_RNO[13]  (.A(\state[1]_net_1 ), 
        .B(\dout[13] ), .Y(N_689_i));
    SLE \pcm_right[4]  (.D(\pcm_right_RNO[4]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[4]));
    SLE \left[21]  (.D(\dout[21] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[21]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \pcm_left_RNO[28]  (.A(\state[1]_net_1 ), 
        .B(use_dsd), .C(\left[28]_net_1 ), .Y(\pcm_left_RNO[28]_net_1 )
        );
    SLE \pcm_right[17]  (.D(N_949_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[17]));
    SLE \pcm_right[7]  (.D(N_749_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[7]));
    SLE \pcm_left[16]  (.D(\pcm_left_RNO[16]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_left[16]));
    SLE \pcm_left[4]  (.D(\pcm_left_RNO[4]_net_1 ), .CLK(mclk_1), .EN(
        un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(source_left[4])
        );
    CFG4 #( .INIT(16'h3C38) )  flag_ldmx (.A(\state[1]_net_1 ), .B(
        flag_en_net_1), .C(flag_net_1), .D(\state[0]_net_1 ), .Y(
        flag_ldmx_net_1));
    SLE \pcm_left[21]  (.D(N_1149_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[21]));
    CFG2 #( .INIT(4'h2) )  n_k20 (.A(in_bck_1), .B(old_bck_net_1), .Y(
        N_162));
    SLE \left[3]  (.D(\dout[3] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \pcm_left_RNO[9]  (.A(\state[1]_net_1 ), .B(
        \left[9]_net_1 ), .Y(N_989_i));
    SLE \pcm_right[13]  (.D(N_689_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_right[13]));
    CFG3 #( .INIT(8'h48) )  k_n1 (.A(\k[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(\k[1]_net_1 ), .Y(k_n1_net_1));
    sync_logic_1s usync100 (.un1_ctrl(un1_ctrl_net_1), 
        .sdctrl_start_i2s(sdctrl_start_i2s), .sdclk_n_1(sdclk_n_1), 
        .mclk_1(mclk_1), .N_4047_i(N_4047_i));
    SLE \pcm_right[12]  (.D(\pcm_right_RNO[12]_net_1 ), .CLK(mclk_1), 
        .EN(un1_state_6_i), .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        source_right[12]));
    SLE \pcm_left[23]  (.D(N_1129_i), .CLK(mclk_1), .EN(un1_state_6_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(source_left[23]));
    CFG3 #( .INIT(8'h60) )  k_n3 (.A(k_c2_net_1), .B(\k[3]_net_1 ), .C(
        \state[1]_net_1 ), .Y(k_n3_net_1));
    SLE sound_card_start (.D(N_3820_i), .CLK(mclk_1), .EN(N_3822_i), 
        .ALn(N_4047_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(i2s_start));
    SLE \left[10]  (.D(\dout[10] ), .CLK(mclk_1), .EN(
        un1_state_7_i_a3_2_net_1), .ALn(N_4047_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \left[10]_net_1 ));
    
endmodule


module pcm_tx(
       source_right,
       source_left,
       reset_n_i_1,
       start_pcm_tx,
       reset_n_i_0_RNIOUJE,
       olrck2,
       odata2,
       in_bck_1,
       reset_n_i_i
    );
input  [31:0] source_right;
input  [31:0] source_left;
output reset_n_i_1;
input  start_pcm_tx;
input  reset_n_i_0_RNIOUJE;
output olrck2;
output odata2;
input  in_bck_1;
input  reset_n_i_i;

    wire \i[0]_net_1 , \i_s[0] , \t1[63]_net_1 , VCC_net_1, 
        \t1_4[63]_net_1 , GND_net_1, \t1[48]_net_1 , \t1_4[48]_net_1 , 
        \t1[49]_net_1 , \t1_4[49]_net_1 , \t1[50]_net_1 , 
        \t1_4_i_m2[50]_net_1 , \t1[51]_net_1 , \t1_4[51]_net_1 , 
        \t1[52]_net_1 , \t1_4_i_m2[52]_net_1 , \t1[53]_net_1 , 
        \t1_4[53]_net_1 , \t1[54]_net_1 , \t1_4_i_m2[54]_net_1 , 
        \t1[55]_net_1 , \t1_4[55]_net_1 , \t1[56]_net_1 , 
        \t1_4[56]_net_1 , \t1[57]_net_1 , \t1_4[57]_net_1 , 
        \t1[58]_net_1 , \t1_4[58]_net_1 , \t1[59]_net_1 , 
        \t1_4[59]_net_1 , \t1[60]_net_1 , \t1_4[60]_net_1 , 
        \t1[61]_net_1 , \t1_4[61]_net_1 , \t1[62]_net_1 , 
        \t1_4[62]_net_1 , \t1[33]_net_1 , \t1_4[33]_net_1 , 
        \t1[34]_net_1 , \t1_4[34]_net_1 , \t1[35]_net_1 , 
        \t1_4[35]_net_1 , \t1[36]_net_1 , \t1_4[36]_net_1 , 
        \t1[37]_net_1 , \t1_4[37]_net_1 , \t1[38]_net_1 , 
        \t1_4[38]_net_1 , \t1[39]_net_1 , \t1_4[39]_net_1 , 
        \t1[40]_net_1 , \t1_4[40]_net_1 , \t1[41]_net_1 , 
        \t1_4[41]_net_1 , \t1[42]_net_1 , \t1_4[42]_net_1 , 
        \t1[43]_net_1 , \t1_4[43]_net_1 , \t1[44]_net_1 , 
        \t1_4[44]_net_1 , \t1[45]_net_1 , \t1_4[45]_net_1 , 
        \t1[46]_net_1 , \t1_4[46]_net_1 , \t1[47]_net_1 , 
        \t1_4[47]_net_1 , \t1[18]_net_1 , \t1_4_i_m2[18]_net_1 , 
        \t1[19]_net_1 , \t1_4[19]_net_1 , \t1[20]_net_1 , 
        \t1_4[20]_net_1 , \t1[21]_net_1 , \t1_4[21]_net_1 , 
        \t1[22]_net_1 , \t1_4_i_m2[22]_net_1 , \t1[23]_net_1 , 
        \t1_4[23]_net_1 , \t1[24]_net_1 , \t1_4[24]_net_1 , 
        \t1[25]_net_1 , \t1_4[25]_net_1 , \t1[26]_net_1 , 
        \t1_4[26]_net_1 , \t1[27]_net_1 , \t1_4[27]_net_1 , 
        \t1[28]_net_1 , \t1_4[28]_net_1 , \t1[29]_net_1 , 
        \t1_4[29]_net_1 , \t1[30]_net_1 , \t1_4[30]_net_1 , 
        \t1[31]_net_1 , \t1_4[31]_net_1 , \t1[32]_net_1 , 
        \t1_4[32]_net_1 , \t1[3]_net_1 , \t1_4[3]_net_1 , 
        \t1[4]_net_1 , \t1_4[4]_net_1 , \t1[5]_net_1 , \t1_4[5]_net_1 , 
        \t1[6]_net_1 , \t1_4[6]_net_1 , \t1[7]_net_1 , \t1_4[7]_net_1 , 
        \t1[8]_net_1 , \t1_4[8]_net_1 , \t1[9]_net_1 , \t1_4[9]_net_1 , 
        \t1[10]_net_1 , \t1_4_i_m2[10]_net_1 , \t1[11]_net_1 , 
        \t1_4[11]_net_1 , \t1[12]_net_1 , \t1_4[12]_net_1 , 
        \t1[13]_net_1 , \t1_4[13]_net_1 , \t1[14]_net_1 , 
        \t1_4[14]_net_1 , \t1[15]_net_1 , \t1_4[15]_net_1 , 
        \t1[16]_net_1 , \t1_4[16]_net_1 , \t1[17]_net_1 , 
        \t1_4[17]_net_1 , \t1[0]_net_1 , \t1_4[0]_net_1 , 
        \t1[1]_net_1 , \t1_4[1]_net_1 , \t1[2]_net_1 , \t1_4[2]_net_1 , 
        \i[1]_net_1 , \i_s[1] , \i[2]_net_1 , \i_s[2] , \i[3]_net_1 , 
        \i_s[3] , \i[4]_net_1 , \i_s[4] , \i_s[5]_net_1 , i_s_414_FCO, 
        \i_cry[1]_net_1 , \i_cry[2]_net_1 , \i_cry[3]_net_1 , 
        \i_cry[4]_net_1 , t19_3_net_1, t19_net_1;
    
    SLE \t1[44]  (.D(\t1_4[44]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[44]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[51]  (.A(t19_net_1), .B(
        \t1[50]_net_1 ), .C(source_left[19]), .Y(\t1_4[51]_net_1 ));
    SLE \t1[0]  (.D(\t1_4[0]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[0]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[30]  (.A(t19_net_1), .B(
        \t1[29]_net_1 ), .C(source_right[30]), .Y(\t1_4[30]_net_1 ));
    SLE \t1[58]  (.D(\t1_4[58]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[58]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[25]  (.A(t19_net_1), .B(
        \t1[24]_net_1 ), .C(source_right[25]), .Y(\t1_4[25]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[61]  (.A(t19_net_1), .B(
        \t1[60]_net_1 ), .C(source_left[29]), .Y(\t1_4[61]_net_1 ));
    SLE \t1[4]  (.D(\t1_4[4]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[4]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[40]  (.A(t19_net_1), .B(
        \t1[39]_net_1 ), .C(source_left[8]), .Y(\t1_4[40]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[4]  (.A(t19_net_1), .B(\t1[3]_net_1 )
        , .C(source_right[4]), .Y(\t1_4[4]_net_1 ));
    SLE \t1[10]  (.D(\t1_4_i_m2[10]_net_1 ), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t1[10]_net_1 ));
    SLE \i[0]  (.D(\i_s[0] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[16]  (.A(t19_net_1), .B(
        \t1[15]_net_1 ), .C(source_right[16]), .Y(\t1_4[16]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_s[5]  (.A(VCC_net_1), .B(olrck2), 
        .C(GND_net_1), .D(GND_net_1), .FCI(\i_cry[4]_net_1 ), .S(
        \i_s[5]_net_1 ), .Y(), .FCO());
    SLE \t1[31]  (.D(\t1_4[31]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[31]_net_1 ));
    SLE \t1[27]  (.D(\t1_4[27]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[27]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[19]  (.A(t19_net_1), .B(
        \t1[18]_net_1 ), .C(source_right[19]), .Y(\t1_4[19]_net_1 ));
    SLE \t1[14]  (.D(\t1_4[14]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[14]_net_1 ));
    SLE \t1[42]  (.D(\t1_4[42]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[42]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[38]  (.A(t19_net_1), .B(
        \t1[37]_net_1 ), .C(source_left[6]), .Y(\t1_4[38]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[17]  (.A(t19_net_1), .B(
        \t1[16]_net_1 ), .C(source_right[17]), .Y(\t1_4[17]_net_1 ));
    SLE \t1[57]  (.D(\t1_4[57]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[57]_net_1 ));
    SLE \t1[63]  (.D(\t1_4[63]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[63]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[48]  (.A(t19_net_1), .B(
        \t1[47]_net_1 ), .C(source_left[16]), .Y(\t1_4[48]_net_1 ));
    CFG3 #( .INIT(8'h80) )  t19 (.A(t19_3_net_1), .B(\i[3]_net_1 ), .C(
        olrck2), .Y(t19_net_1));
    SLE \t1[7]  (.D(\t1_4[7]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[7]_net_1 ));
    SLE \t1[39]  (.D(\t1_4[39]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[39]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \t1[26]  (.D(\t1_4[26]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[26]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[33]  (.A(t19_net_1), .B(
        \t1[32]_net_1 ), .C(source_left[1]), .Y(\t1_4[33]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[24]  (.A(t19_net_1), .B(
        \t1[23]_net_1 ), .C(source_right[24]), .Y(\t1_4[24]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[56]  (.A(t19_net_1), .B(
        \t1[55]_net_1 ), .C(source_left[24]), .Y(\t1_4[56]_net_1 ));
    SLE \t1[45]  (.D(\t1_4[45]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[45]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[59]  (.A(t19_net_1), .B(
        \t1[58]_net_1 ), .C(source_left[27]), .Y(\t1_4[59]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \i_RNO[0]  (.A(\i[0]_net_1 ), .Y(\i_s[0] ));
    SLE d1 (.D(\t1[63]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(odata2));
    CFG3 #( .INIT(8'hE4) )  \t1_4[43]  (.A(t19_net_1), .B(
        \t1[42]_net_1 ), .C(source_left[11]), .Y(\t1_4[43]_net_1 ));
    SLE \t1[60]  (.D(\t1_4[60]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[60]_net_1 ));
    SLE \t1[56]  (.D(\t1_4[56]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[56]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[6]  (.A(t19_net_1), .B(\t1[5]_net_1 )
        , .C(source_right[6]), .Y(\t1_4[6]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[35]  (.A(t19_net_1), .B(
        \t1[34]_net_1 ), .C(source_left[3]), .Y(\t1_4[35]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[57]  (.A(t19_net_1), .B(
        \t1[56]_net_1 ), .C(source_left[25]), .Y(\t1_4[57]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4_i_m2[50]  (.A(t19_net_1), .B(
        \t1[49]_net_1 ), .C(source_left[18]), .Y(\t1_4_i_m2[50]_net_1 )
        );
    SLE \t1[23]  (.D(\t1_4[23]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[23]_net_1 ));
    SLE \t1[12]  (.D(\t1_4[12]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[12]_net_1 ));
    SLE \t1[38]  (.D(\t1_4[38]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[38]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[45]  (.A(t19_net_1), .B(
        \t1[44]_net_1 ), .C(source_left[13]), .Y(\t1_4[45]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[21]  (.A(t19_net_1), .B(
        \t1[20]_net_1 ), .C(source_right[21]), .Y(\t1_4[21]_net_1 ));
    SLE \t1[53]  (.D(\t1_4[53]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[53]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4_i_m2[52]  (.A(t19_net_1), .B(
        \t1[51]_net_1 ), .C(source_left[20]), .Y(\t1_4_i_m2[52]_net_1 )
        );
    SLE \t1[3]  (.D(\t1_4[3]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[3]_net_1 ));
    SLE \t1[20]  (.D(\t1_4[20]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[20]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[12]  (.A(t19_net_1), .B(
        \t1[11]_net_1 ), .C(source_right[12]), .Y(\t1_4[12]_net_1 ));
    SLE \t1[15]  (.D(\t1_4[15]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[15]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \t1[50]  (.D(\t1_4_i_m2[50]_net_1 ), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t1[50]_net_1 ));
    SLE \t1[37]  (.D(\t1_4[37]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[37]_net_1 ));
    SLE \t1[24]  (.D(\t1_4[24]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[24]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[34]  (.A(t19_net_1), .B(
        \t1[33]_net_1 ), .C(source_left[2]), .Y(\t1_4[34]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[7]  (.A(t19_net_1), .B(\t1[6]_net_1 )
        , .C(source_right[7]), .Y(\t1_4[7]_net_1 ));
    SLE \t1[54]  (.D(\t1_4_i_m2[54]_net_1 ), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t1[54]_net_1 ));
    SLE \t1[62]  (.D(\t1_4[62]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[62]_net_1 ));
    SLE \t1[41]  (.D(\t1_4[41]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[41]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[44]  (.A(t19_net_1), .B(
        \t1[43]_net_1 ), .C(source_left[12]), .Y(\t1_4[44]_net_1 ));
    SLE \t1[6]  (.D(\t1_4[6]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[6]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[62]  (.A(t19_net_1), .B(
        \t1[61]_net_1 ), .C(source_left[30]), .Y(\t1_4[62]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[26]  (.A(t19_net_1), .B(
        \t1[25]_net_1 ), .C(source_right[26]), .Y(\t1_4[26]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  t19_3 (.A(\i[4]_net_1 ), .B(
        \i[2]_net_1 ), .C(\i[1]_net_1 ), .D(\i[0]_net_1 ), .Y(
        t19_3_net_1));
    CFG3 #( .INIT(8'hE4) )  \t1_4[29]  (.A(t19_net_1), .B(
        \t1[28]_net_1 ), .C(source_right[29]), .Y(\t1_4[29]_net_1 ));
    SLE \t1[36]  (.D(\t1_4[36]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[36]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[31]  (.A(t19_net_1), .B(
        \t1[30]_net_1 ), .C(source_right[31]), .Y(\t1_4[31]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[27]  (.A(t19_net_1), .B(
        \t1[26]_net_1 ), .C(source_right[27]), .Y(\t1_4[27]_net_1 ));
    SLE \t1[2]  (.D(\t1_4[2]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[2]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[41]  (.A(t19_net_1), .B(
        \t1[40]_net_1 ), .C(source_left[9]), .Y(\t1_4[41]_net_1 ));
    SLE \t1[49]  (.D(\t1_4[49]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[49]_net_1 ));
    SLE \t1[22]  (.D(\t1_4_i_m2[22]_net_1 ), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t1[22]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4_i_m2[10]  (.A(t19_net_1), .B(
        \t1[9]_net_1 ), .C(source_right[10]), .Y(\t1_4_i_m2[10]_net_1 )
        );
    SLE \t1[33]  (.D(\t1_4[33]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[33]_net_1 ));
    SLE \i[2]  (.D(\i_s[2] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    SLE \t1[11]  (.D(\t1_4[11]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[11]_net_1 ));
    SLE \t1[52]  (.D(\t1_4_i_m2[52]_net_1 ), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t1[52]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[60]  (.A(t19_net_1), .B(
        \t1[59]_net_1 ), .C(source_left[28]), .Y(\t1_4[60]_net_1 ));
    SLE \t1[48]  (.D(\t1_4[48]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[48]_net_1 ));
    SLE \t1[25]  (.D(\t1_4[25]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[25]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4_i_m2[54]  (.A(t19_net_1), .B(
        \t1[53]_net_1 ), .C(source_left[22]), .Y(\t1_4_i_m2[54]_net_1 )
        );
    SLE \t1[30]  (.D(\t1_4[30]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[30]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[13]  (.A(t19_net_1), .B(
        \t1[12]_net_1 ), .C(source_right[13]), .Y(\t1_4[13]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(i_s_414_FCO), 
        .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[4]  (.D(\i_s[4] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    SLE \t1[55]  (.D(\t1_4[55]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[55]_net_1 ));
    SLE \t1[19]  (.D(\t1_4[19]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[19]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[15]  (.A(t19_net_1), .B(
        \t1[14]_net_1 ), .C(source_right[15]), .Y(\t1_4[15]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[58]  (.A(t19_net_1), .B(
        \t1[57]_net_1 ), .C(source_left[26]), .Y(\t1_4[58]_net_1 ));
    CFG2 #( .INIT(4'h4) )  reset_n_i (.A(reset_n_i_0_RNIOUJE), .B(
        start_pcm_tx), .Y(reset_n_i_1));
    SLE \t1[34]  (.D(\t1_4[34]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[34]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[36]  (.A(t19_net_1), .B(
        \t1[35]_net_1 ), .C(source_left[4]), .Y(\t1_4[36]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[39]  (.A(t19_net_1), .B(
        \t1[38]_net_1 ), .C(source_left[7]), .Y(\t1_4[39]_net_1 ));
    SLE \t1[5]  (.D(\t1_4[5]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[5]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[46]  (.A(t19_net_1), .B(
        \t1[45]_net_1 ), .C(source_left[14]), .Y(\t1_4[46]_net_1 ));
    SLE \t1[47]  (.D(\t1_4[47]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[47]_net_1 ));
    SLE \t1[18]  (.D(\t1_4_i_m2[18]_net_1 ), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t1[18]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[53]  (.A(t19_net_1), .B(
        \t1[52]_net_1 ), .C(source_left[21]), .Y(\t1_4[53]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[49]  (.A(t19_net_1), .B(
        \t1[48]_net_1 ), .C(source_left[17]), .Y(\t1_4[49]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[37]  (.A(t19_net_1), .B(
        \t1[36]_net_1 ), .C(source_left[5]), .Y(\t1_4[37]_net_1 ));
    SLE \t1[61]  (.D(\t1_4[61]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[61]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[63]  (.A(t19_net_1), .B(
        \t1[62]_net_1 ), .C(source_left[31]), .Y(\t1_4[63]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[47]  (.A(t19_net_1), .B(
        \t1[46]_net_1 ), .C(source_left[15]), .Y(\t1_4[47]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[55]  (.A(t19_net_1), .B(
        \t1[54]_net_1 ), .C(source_left[23]), .Y(\t1_4[55]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[5]  (.A(t19_net_1), .B(\t1[4]_net_1 )
        , .C(source_right[5]), .Y(\t1_4[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    SLE \i[5]  (.D(\i_s[5]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(olrck2));
    CFG3 #( .INIT(8'hE4) )  \t1_4[20]  (.A(t19_net_1), .B(
        \t1[19]_net_1 ), .C(source_right[20]), .Y(\t1_4[20]_net_1 ));
    SLE \t1[32]  (.D(\t1_4[32]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[32]_net_1 ));
    SLE \t1[46]  (.D(\t1_4[46]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[46]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4_i_m2[18]  (.A(t19_net_1), .B(
        \t1[17]_net_1 ), .C(source_right[18]), .Y(
        \t1_4_i_m2[18]_net_1 ));
    SLE \t1[21]  (.D(\t1_4[21]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[21]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[14]  (.A(t19_net_1), .B(
        \t1[13]_net_1 ), .C(source_right[14]), .Y(\t1_4[14]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[8]  (.A(t19_net_1), .B(\t1[7]_net_1 )
        , .C(source_right[8]), .Y(\t1_4[8]_net_1 ));
    SLE \t1[17]  (.D(\t1_4[17]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[17]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[9]  (.A(t19_net_1), .B(\t1[8]_net_1 )
        , .C(source_right[9]), .Y(\t1_4[9]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[2]  (.A(t19_net_1), .B(\t1[1]_net_1 )
        , .C(source_right[2]), .Y(\t1_4[2]_net_1 ));
    SLE \t1[51]  (.D(\t1_4[51]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[51]_net_1 ));
    SLE \t1[43]  (.D(\t1_4[43]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[43]_net_1 ));
    SLE \i[3]  (.D(\i_s[3] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    SLE \t1[35]  (.D(\t1_4[35]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[35]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[11]  (.A(t19_net_1), .B(
        \t1[10]_net_1 ), .C(source_right[11]), .Y(\t1_4[11]_net_1 ));
    SLE \t1[29]  (.D(\t1_4[29]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[29]_net_1 ));
    SLE \i[1]  (.D(\i_s[1] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4_i_m2[22]  (.A(t19_net_1), .B(
        \t1[21]_net_1 ), .C(source_right[22]), .Y(
        \t1_4_i_m2[22]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[32]  (.A(t19_net_1), .B(
        \t1[31]_net_1 ), .C(source_left[0]), .Y(\t1_4[32]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[28]  (.A(t19_net_1), .B(
        \t1[27]_net_1 ), .C(source_right[28]), .Y(\t1_4[28]_net_1 ));
    SLE \t1[16]  (.D(\t1_4[16]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[16]_net_1 ));
    SLE \t1[40]  (.D(\t1_4[40]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[40]_net_1 ));
    SLE \t1[9]  (.D(\t1_4[9]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[9]_net_1 ));
    SLE \t1[59]  (.D(\t1_4[59]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[59]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[42]  (.A(t19_net_1), .B(
        \t1[41]_net_1 ), .C(source_left[10]), .Y(\t1_4[42]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[3]  (.A(t19_net_1), .B(\t1[2]_net_1 )
        , .C(source_right[3]), .Y(\t1_4[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  i_s_414 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(i_s_414_FCO));
    CFG4 #( .INIT(16'h8000) )  \t1_4[0]  (.A(olrck2), .B(\i[3]_net_1 ), 
        .C(t19_3_net_1), .D(source_right[0]), .Y(\t1_4[0]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[1]  (.A(t19_net_1), .B(\t1[0]_net_1 )
        , .C(source_right[1]), .Y(\t1_4[1]_net_1 ));
    SLE \t1[8]  (.D(\t1_4[8]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[8]_net_1 ));
    SLE \t1[28]  (.D(\t1_4[28]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[28]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \t1_4[23]  (.A(t19_net_1), .B(
        \t1[22]_net_1 ), .C(source_right[23]), .Y(\t1_4[23]_net_1 ));
    SLE \t1[1]  (.D(\t1_4[1]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[1]_net_1 ));
    SLE \t1[13]  (.D(\t1_4[13]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[13]_net_1 ));
    
endmodule


module dsd_tx(
       source_left,
       source_right,
       reset_n_i_0,
       start_dsd_tx,
       reset_n_i_0_RNIOUJE,
       odata1,
       olrck1,
       dsd_clk_1,
       reset_n_i_i
    );
input  [31:0] source_left;
input  [31:0] source_right;
output reset_n_i_0;
input  start_dsd_tx;
input  reset_n_i_0_RNIOUJE;
output odata1;
output olrck1;
input  dsd_clk_1;
input  reset_n_i_i;

    wire \i[0]_net_1 , \i_i[0] , VCC_net_1, GND_net_1, \i[1]_net_1 , 
        N_36_i, \i[2]_net_1 , N_37_i_i, \i[3]_net_1 , N_38_i_i, 
        \i[4]_net_1 , N_39_i_i, \t1[21]_net_1 , \t1_4[21]_net_1 , 
        \t1[22]_net_1 , \t1_4[22]_net_1 , \t1[23]_net_1 , 
        \t1_4[23]_net_1 , \t1[24]_net_1 , \t1_4[24]_net_1 , 
        \t1[25]_net_1 , \t1_4[25]_net_1 , \t1[26]_net_1 , 
        \t1_4[26]_net_1 , \t1[27]_net_1 , \t1_4[27]_net_1 , 
        \t1[28]_net_1 , \t1_4[28]_net_1 , \t1[29]_net_1 , 
        \t1_4[29]_net_1 , \t1[30]_net_1 , \t1_4[30]_net_1 , 
        \t1_4[31]_net_1 , \t1[6]_net_1 , \t1_4[6]_net_1 , 
        \t1[7]_net_1 , \t1_4[7]_net_1 , \t1[8]_net_1 , \t1_4[8]_net_1 , 
        \t1[9]_net_1 , \t1_4[9]_net_1 , \t1[10]_net_1 , 
        \t1_4[10]_net_1 , \t1[11]_net_1 , \t1_4[11]_net_1 , 
        \t1[12]_net_1 , \t1_4[12]_net_1 , \t1[13]_net_1 , 
        \t1_4[13]_net_1 , \t1[14]_net_1 , \t1_4[14]_net_1 , 
        \t1[15]_net_1 , \t1_4[15]_net_1 , \t1[16]_net_1 , 
        \t1_4[16]_net_1 , \t1[17]_net_1 , \t1_4[17]_net_1 , 
        \t1[18]_net_1 , \t1_4[18]_net_1 , \t1[19]_net_1 , 
        \t1_4[19]_net_1 , \t1[20]_net_1 , \t1_4[20]_net_1 , 
        \t2[23]_net_1 , \t2_4[23]_net_1 , \t2[24]_net_1 , 
        \t2_4[24]_net_1 , \t2[25]_net_1 , \t2_4[25]_net_1 , 
        \t2[26]_net_1 , \t2_4[26]_net_1 , \t2[27]_net_1 , 
        \t2_4[27]_net_1 , \t2[28]_net_1 , \t2_4[28]_net_1 , 
        \t2[29]_net_1 , \t2_4[29]_net_1 , \t2[30]_net_1 , 
        \t2_4[30]_net_1 , \t2_4[31]_net_1 , \t1[0]_net_1 , 
        \t1_4[0]_net_1 , \t1[1]_net_1 , \t1_4[1]_net_1 , \t1[2]_net_1 , 
        \t1_4[2]_net_1 , \t1[3]_net_1 , \t1_4[3]_net_1 , \t1[4]_net_1 , 
        \t1_4[4]_net_1 , \t1[5]_net_1 , \t1_4[5]_net_1 , \t2[8]_net_1 , 
        \t2_4[8]_net_1 , \t2[9]_net_1 , \t2_4[9]_net_1 , 
        \t2[10]_net_1 , \t2_4_i_m2[10]_net_1 , \t2[11]_net_1 , 
        \t2_4[11]_net_1 , \t2[12]_net_1 , \t2_4[12]_net_1 , 
        \t2[13]_net_1 , \t2_4[13]_net_1 , \t2[14]_net_1 , 
        \t2_4[14]_net_1 , \t2[15]_net_1 , \t2_4[15]_net_1 , 
        \t2[16]_net_1 , \t2_4[16]_net_1 , \t2[17]_net_1 , 
        \t2_4[17]_net_1 , \t2[18]_net_1 , \t2_4_i_m2[18]_net_1 , 
        \t2[19]_net_1 , \t2_4[19]_net_1 , \t2[20]_net_1 , 
        \t2_4[20]_net_1 , \t2[21]_net_1 , \t2_4[21]_net_1 , 
        \t2[22]_net_1 , \t2_4_i_m2[22]_net_1 , \t2[0]_net_1 , 
        \t2_4[0]_net_1 , \t2[1]_net_1 , \t2_4[1]_net_1 , \t2[2]_net_1 , 
        \t2_4[2]_net_1 , \t2[3]_net_1 , \t2_4[3]_net_1 , \t2[4]_net_1 , 
        \t2_4[4]_net_1 , \t2[5]_net_1 , \t2_4[5]_net_1 , \t2[6]_net_1 , 
        \t2_4[6]_net_1 , \t2[7]_net_1 , \t2_4[7]_net_1 , N_3911;
    
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[7]  (.A(source_right[7]), .B(
        \t2[6]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[7]_net_1 ));
    CFG3 #( .INIT(8'h6A) )  \i_RNO[2]  (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(\i[0]_net_1 ), .Y(N_37_i_i));
    SLE \t1[0]  (.D(\t1_4[0]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[0]_net_1 ));
    SLE \t2[10]  (.D(\t2_4_i_m2[10]_net_1 ), .CLK(dsd_clk_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t2[10]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[30]  (.A(source_left[30]), .B(
        \t1[29]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[30]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[30]  (.A(source_right[30]), .B(
        \t2[29]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[30]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[25]  (.A(source_left[25]), .B(
        \t1[24]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[25]_net_1 ));
    SLE \t1[4]  (.D(\t1_4[4]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[4]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[24]  (.A(source_right[24]), .B(
        \t2[23]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[24]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[8]  (.A(source_right[8]), .B(
        \t2[7]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[8]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[12]  (.A(source_right[12]), .B(
        \t2[11]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[12]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[4]  (.A(source_left[4]), .B(
        \t1[3]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[4]_net_1 ));
    SLE \t2[7]  (.D(\t2_4[7]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[7]_net_1 ));
    SLE \t2[3]  (.D(\t2_4[3]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[3]_net_1 ));
    SLE \t1[10]  (.D(\t1_4[10]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[10]_net_1 ));
    SLE \i[0]  (.D(\i_i[0] ), .CLK(dsd_clk_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    SLE \t2[14]  (.D(\t2_4[14]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[14]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[1]  (.A(source_right[1]), .B(
        \t2[0]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[1]_net_1 ));
    CFG4 #( .INIT(16'h6AAA) )  \i_RNO[3]  (.A(\i[3]_net_1 ), .B(
        \i[2]_net_1 ), .C(\i[1]_net_1 ), .D(\i[0]_net_1 ), .Y(N_38_i_i)
        );
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[16]  (.A(source_left[16]), .B(
        \t1[15]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[16]_net_1 ));
    SLE \t1[31]  (.D(\t1_4[31]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(olrck1));
    SLE \t1[27]  (.D(\t1_4[27]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[27]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[19]  (.A(source_left[19]), .B(
        \t1[18]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[19]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[21]  (.A(source_right[21]), .B(
        \t2[20]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[21]_net_1 ));
    CFG2 #( .INIT(4'h9) )  \i_RNO[4]  (.A(N_3911), .B(\i[4]_net_1 ), 
        .Y(N_39_i_i));
    SLE \t2[22]  (.D(\t2_4_i_m2[22]_net_1 ), .CLK(dsd_clk_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t2[22]_net_1 ));
    SLE \t1[14]  (.D(\t1_4[14]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[14]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[17]  (.A(source_left[17]), .B(
        \t1[16]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[17]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[6]  (.A(source_right[6]), .B(
        \t2[5]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[6]_net_1 ));
    SLE \t1[7]  (.D(\t1_4[7]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[7]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \t1[26]  (.D(\t1_4[26]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[26]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[24]  (.A(source_left[24]), .B(
        \t1[23]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[24]_net_1 ));
    SLE \t2[25]  (.D(\t2_4[25]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[25]_net_1 ));
    SLE \t2[12]  (.D(\t2_4[12]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[12]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \i_RNO[0]  (.A(\i[0]_net_1 ), .Y(\i_i[0] ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[6]  (.A(source_left[6]), .B(
        \t1[5]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[6]_net_1 ));
    SLE \t1[23]  (.D(\t1_4[23]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[23]_net_1 ));
    SLE \t1[12]  (.D(\t1_4[12]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[12]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[21]  (.A(source_left[21]), .B(
        \t1[20]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[21]_net_1 ));
    SLE \t2[15]  (.D(\t2_4[15]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[15]_net_1 ));
    SLE \t2[0]  (.D(\t2_4[0]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[0]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[26]  (.A(source_right[26]), .B(
        \t2[25]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[26]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[4]  (.A(source_right[4]), .B(
        \t2[3]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[4]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[29]  (.A(source_right[29]), .B(
        \t2[28]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[29]_net_1 ));
    SLE \t1[3]  (.D(\t1_4[3]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[3]_net_1 ));
    SLE \t1[20]  (.D(\t1_4[20]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[20]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4_i_m2[22]  (.A(source_right[22]), 
        .B(\t2[21]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4_i_m2[22]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[13]  (.A(source_right[13]), .B(
        \t2[12]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[13]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[12]  (.A(source_left[12]), .B(
        \t1[11]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[12]_net_1 ));
    SLE \t1[15]  (.D(\t1_4[15]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[15]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[27]  (.A(source_right[27]), .B(
        \t2[26]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[27]_net_1 ));
    SLE \t2[31]  (.D(\t2_4[31]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(odata1));
    SLE \t2[2]  (.D(\t2_4[2]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[2]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \t2_4[0]  (.A(source_right[0]), .B(
        \i[4]_net_1 ), .C(N_3911), .Y(\t2_4[0]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[15]  (.A(source_right[15]), .B(
        \t2[14]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[15]_net_1 ));
    SLE \t2[6]  (.D(\t2_4[6]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[6]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[2]  (.A(source_right[2]), .B(
        \t2[1]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[2]_net_1 ));
    SLE \t1[24]  (.D(\t1_4[24]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[24]_net_1 ));
    SLE \t2[21]  (.D(\t2_4[21]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[21]_net_1 ));
    SLE \t2[9]  (.D(\t2_4[9]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[9]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[7]  (.A(source_left[7]), .B(
        \t1[6]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[7]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[10]  (.A(source_left[10]), .B(
        \t1[9]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[10]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  t19_0_o4 (.A(\i[3]_net_1 ), .B(
        \i[2]_net_1 ), .C(\i[1]_net_1 ), .D(\i[0]_net_1 ), .Y(N_3911));
    SLE \t1[6]  (.D(\t1_4[6]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[6]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[26]  (.A(source_left[26]), .B(
        \t1[25]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[26]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[29]  (.A(source_left[29]), .B(
        \t1[28]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[29]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[31]  (.A(source_left[31]), .B(
        \t1[30]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[31]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[31]  (.A(source_right[31]), .B(
        \t2[30]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[31]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[27]  (.A(source_left[27]), .B(
        \t1[26]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[27]_net_1 ));
    SLE \t1[2]  (.D(\t1_4[2]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[2]_net_1 ));
    SLE \t2[29]  (.D(\t2_4[29]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[29]_net_1 ));
    SLE \t2[11]  (.D(\t2_4[11]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[11]_net_1 ));
    SLE \t1[22]  (.D(\t1_4[22]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[22]_net_1 ));
    SLE \i[2]  (.D(N_37_i_i), .CLK(dsd_clk_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[14]  (.A(source_right[14]), .B(
        \t2[13]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[14]_net_1 ));
    SLE \t2[8]  (.D(\t2_4[8]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[8]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[18]  (.A(source_left[18]), .B(
        \t1[17]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[18]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[5]  (.A(source_right[5]), .B(
        \t2[4]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[5]_net_1 ));
    SLE \t1[11]  (.D(\t1_4[11]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[11]_net_1 ));
    SLE \t2[28]  (.D(\t2_4[28]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[28]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4_i_m2[18]  (.A(source_right[18]), 
        .B(\t2[17]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4_i_m2[18]_net_1 ));
    SLE \t1[25]  (.D(\t1_4[25]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[25]_net_1 ));
    SLE \t2[19]  (.D(\t2_4[19]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[19]_net_1 ));
    SLE \t1[30]  (.D(\t1_4[30]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[30]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[13]  (.A(source_left[13]), .B(
        \t1[12]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[13]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[11]  (.A(source_right[11]), .B(
        \t2[10]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[11]_net_1 ));
    SLE \i[4]  (.D(N_39_i_i), .CLK(dsd_clk_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    SLE \t1[19]  (.D(\t1_4[19]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[19]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[20]  (.A(source_right[20]), .B(
        \t2[19]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[20]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[15]  (.A(source_left[15]), .B(
        \t1[14]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[15]_net_1 ));
    CFG2 #( .INIT(4'h4) )  reset_n_i (.A(reset_n_i_0_RNIOUJE), .B(
        start_dsd_tx), .Y(reset_n_i_0));
    SLE \t2[18]  (.D(\t2_4_i_m2[18]_net_1 ), .CLK(dsd_clk_1), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\t2[18]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[22]  (.A(source_left[22]), .B(
        \t1[21]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[22]_net_1 ));
    SLE \t2[27]  (.D(\t2_4[27]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[27]_net_1 ));
    SLE \t1[5]  (.D(\t1_4[5]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[5]_net_1 ));
    SLE \t1[18]  (.D(\t1_4[18]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[18]_net_1 ));
    CFG2 #( .INIT(4'h6) )  i_n1_0_x4 (.A(\i[0]_net_1 ), .B(
        \i[1]_net_1 ), .Y(N_36_i));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[28]  (.A(source_right[28]), .B(
        \t2[27]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[28]_net_1 ));
    SLE \t2[5]  (.D(\t2_4[5]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[5]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[5]  (.A(source_left[5]), .B(
        \t1[4]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[5]_net_1 ));
    SLE \t2[1]  (.D(\t2_4[1]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[1]_net_1 ));
    SLE \t2[17]  (.D(\t2_4[17]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[17]_net_1 ));
    SLE \t2[26]  (.D(\t2_4[26]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[26]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[20]  (.A(source_left[20]), .B(
        \t1[19]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[20]_net_1 ));
    SLE \t2[4]  (.D(\t2_4[4]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[4]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[16]  (.A(source_right[16]), .B(
        \t2[15]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[16]_net_1 ));
    SLE \t1[21]  (.D(\t1_4[21]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[21]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[23]  (.A(source_right[23]), .B(
        \t2[22]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[23]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[19]  (.A(source_right[19]), .B(
        \t2[18]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[19]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[14]  (.A(source_left[14]), .B(
        \t1[13]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[14]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[3]  (.A(source_right[3]), .B(
        \t2[2]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[3]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[8]  (.A(source_left[8]), .B(
        \t1[7]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[8]_net_1 ));
    SLE \t1[17]  (.D(\t1_4[17]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[17]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[9]  (.A(source_left[9]), .B(
        \t1[8]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[9]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[2]  (.A(source_left[2]), .B(
        \t1[1]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[2]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[17]  (.A(source_right[17]), .B(
        \t2[16]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[17]_net_1 ));
    SLE \t2[23]  (.D(\t2_4[23]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[23]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[25]  (.A(source_right[25]), .B(
        \t2[24]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[25]_net_1 ));
    SLE \t2[30]  (.D(\t2_4[30]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[30]_net_1 ));
    SLE \i[3]  (.D(N_38_i_i), .CLK(dsd_clk_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    SLE \t2[16]  (.D(\t2_4[16]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[16]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[11]  (.A(source_left[11]), .B(
        \t1[10]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[11]_net_1 ));
    SLE \t1[29]  (.D(\t1_4[29]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[29]_net_1 ));
    SLE \i[1]  (.D(N_36_i), .CLK(dsd_clk_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[28]  (.A(source_left[28]), .B(
        \t1[27]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[28]_net_1 ));
    SLE \t2[20]  (.D(\t2_4[20]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[20]_net_1 ));
    SLE \t1[16]  (.D(\t1_4[16]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[16]_net_1 ));
    SLE \t1[9]  (.D(\t1_4[9]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[9]_net_1 ));
    SLE \t2[13]  (.D(\t2_4[13]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[13]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4_i_m2[10]  (.A(source_right[10]), 
        .B(\t2[9]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4_i_m2[10]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[3]  (.A(source_left[3]), .B(
        \t1[2]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[3]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \t1_4[0]  (.A(source_left[0]), .B(
        \i[4]_net_1 ), .C(N_3911), .Y(\t1_4[0]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[1]  (.A(source_left[1]), .B(
        \t1[0]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[1]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t2_4[9]  (.A(source_right[9]), .B(
        \t2[8]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t2_4[9]_net_1 ));
    SLE \t1[8]  (.D(\t1_4[8]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[8]_net_1 ));
    SLE \t1[28]  (.D(\t1_4[28]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[28]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  \t1_4[23]  (.A(source_left[23]), .B(
        \t1[22]_net_1 ), .C(\i[4]_net_1 ), .D(N_3911), .Y(
        \t1_4[23]_net_1 ));
    SLE \t1[1]  (.D(\t1_4[1]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[1]_net_1 ));
    SLE \t1[13]  (.D(\t1_4[13]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t1[13]_net_1 ));
    SLE \t2[24]  (.D(\t2_4[24]_net_1 ), .CLK(dsd_clk_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\t2[24]_net_1 ));
    
endmodule


module clock_divider(
       dsd138_ctrl,
       bcko,
       N_67,
       bckox4_sn_N_3,
       start_pcm_tx_2,
       dop_start,
       use_dsd,
       i2s_start,
       N_68,
       bckox2,
       clk8,
       clk4,
       mclk_1,
       reset_n_i_i
    );
input  [2:0] dsd138_ctrl;
output bcko;
output N_67;
output bckox4_sn_N_3;
output start_pcm_tx_2;
output dop_start;
input  use_dsd;
input  i2s_start;
output N_68;
output bckox2;
output clk8;
output clk4;
input  mclk_1;
input  reset_n_i_i;

    wire clk32_net_1, clk32_i, clk16_i_i, clk8_i_i, clk4_i_i, clk2_i_i, 
        VCC_net_1, GND_net_1, clk2_net_1, clk16_net_1, 
        bckox2_6_0_0_wmux_0_Y, bckox2_6_0_0_y0, bckox2_6_0_0_co0, N_79, 
        bcko_3_0_0_y0, bcko_3_0_0_co0, bckox2_6_2_net_1, bcko_5_1_0, 
        N_81, bckox2_6_3_net_1;
    
    CFG2 #( .INIT(4'h2) )  bckox4_sn_m2 (.A(dsd138_ctrl[0]), .B(
        dsd138_ctrl[1]), .Y(bckox4_sn_N_3));
    CFG3 #( .INIT(8'h98) )  bckox2_6_2 (.A(dsd138_ctrl[1]), .B(
        dsd138_ctrl[0]), .C(mclk_1), .Y(bckox2_6_2_net_1));
    CFG1 #( .INIT(2'h1) )  clk2_RNO (.A(clk2_net_1), .Y(clk2_i_i));
    ARI1 #( .INIT(20'h0F588) )  bcko_3_0_0_wmux_0 (.A(bcko_3_0_0_y0), 
        .B(dsd138_ctrl[1]), .C(clk8), .D(clk4), .FCI(bcko_3_0_0_co0), 
        .S(), .Y(N_79), .FCO());
    ARI1 #( .INIT(20'h0FA44) )  bcko_3_0_0_wmux (.A(dsd138_ctrl[0]), 
        .B(dsd138_ctrl[1]), .C(clk32_net_1), .D(clk16_net_1), .FCI(
        VCC_net_1), .S(), .Y(bcko_3_0_0_y0), .FCO(bcko_3_0_0_co0));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hC808) )  bckox4_2 (.A(clk2_net_1), .B(
        dsd138_ctrl[1]), .C(dsd138_ctrl[0]), .D(mclk_1), .Y(N_67));
    CFG2 #( .INIT(4'h8) )  dop_start_inst_1 (.A(i2s_start), .B(use_dsd)
        , .Y(dop_start));
    CFG1 #( .INIT(2'h1) )  clk8_RNO (.A(clk8), .Y(clk8_i_i));
    CFG3 #( .INIT(8'hD8) )  bckox2_6_3_RNIONB81 (.A(dsd138_ctrl[2]), 
        .B(bckox2_6_3_net_1), .C(bckox2_6_0_0_wmux_0_Y), .Y(bckox2));
    CFG1 #( .INIT(2'h1) )  clk32_RNO (.A(clk32_net_1), .Y(clk32_i));
    SLE clk32 (.D(clk32_i), .CLK(clk16_net_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(clk32_net_1));
    SLE clk2 (.D(clk2_i_i), .CLK(mclk_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(clk2_net_1));
    CFG3 #( .INIT(8'hB8) )  bckox2_6_3 (.A(clk16_net_1), .B(
        dsd138_ctrl[1]), .C(bckox2_6_2_net_1), .Y(bckox2_6_3_net_1));
    ARI1 #( .INIT(20'h0F588) )  bckox2_6_0_0_wmux_0 (.A(
        bckox2_6_0_0_y0), .B(dsd138_ctrl[1]), .C(clk4), .D(clk2_net_1), 
        .FCI(bckox2_6_0_0_co0), .S(), .Y(bckox2_6_0_0_wmux_0_Y), .FCO()
        );
    CFG3 #( .INIT(8'hD8) )  bcko_6 (.A(dsd138_ctrl[2]), .B(N_81), .C(
        N_79), .Y(bcko));
    CFG1 #( .INIT(2'h1) )  clk4_RNO (.A(clk4), .Y(clk4_i_i));
    SLE clk4_inst_1 (.D(clk4_i_i), .CLK(clk2_net_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(clk4));
    CFG1 #( .INIT(2'h1) )  clk16_RNO (.A(clk16_net_1), .Y(clk16_i_i));
    SLE clk16 (.D(clk16_i_i), .CLK(clk8), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(clk16_net_1));
    CFG3 #( .INIT(8'hC5) )  bcko_5 (.A(bcko_5_1_0), .B(clk32_net_1), 
        .C(dsd138_ctrl[1]), .Y(N_81));
    ARI1 #( .INIT(20'h0FA44) )  bckox2_6_0_0_wmux (.A(dsd138_ctrl[0]), 
        .B(dsd138_ctrl[1]), .C(clk16_net_1), .D(clk8), .FCI(VCC_net_1), 
        .S(), .Y(bckox2_6_0_0_y0), .FCO(bckox2_6_0_0_co0));
    CFG3 #( .INIT(8'h47) )  bcko_5_1 (.A(mclk_1), .B(dsd138_ctrl[0]), 
        .C(clk2_net_1), .Y(bcko_5_1_0));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h2) )  start_pcm_tx_2_inst_1 (.A(i2s_start), .B(
        use_dsd), .Y(start_pcm_tx_2));
    SLE clk8_inst_1 (.D(clk8_i_i), .CLK(clk4), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(clk8));
    CFG2 #( .INIT(4'h6) )  bckox4_sn_m3 (.A(dsd138_ctrl[1]), .B(
        dsd138_ctrl[2]), .Y(N_68));
    
endmodule


module inctrl(
       dsd138_ctrl,
       cnt_0,
       mclk_1,
       dop_start,
       start_pcm_tx_2,
       dop_clock_0,
       spdif_clock_0,
       master_lrck,
       i2s_start,
       use_dsd,
       in_bck_1,
       reset_n_i_i
    );
input  [2:0] dsd138_ctrl;
output cnt_0;
input  mclk_1;
output dop_start;
output start_pcm_tx_2;
output dop_clock_0;
output spdif_clock_0;
output master_lrck;
input  i2s_start;
input  use_dsd;
output in_bck_1;
input  reset_n_i_i;

    wire \cnt[0]_net_1 , \cnt_s[0] , VCC_net_1, GND_net_1, 
        \cnt[1]_net_1 , \cnt_s[1] , \cnt[2]_net_1 , \cnt_s[2] , 
        \cnt[3]_net_1 , \cnt_s[3] , \cnt[4]_net_1 , \cnt_s[4] , 
        \cnt_s[5]_net_1 , cnt_s_415_FCO, \cnt_cry[1]_net_1 , 
        \cnt_cry[2]_net_1 , \cnt_cry[3]_net_1 , \cnt_cry[4]_net_1 , 
        N_68, bckox2, un1_bckox2_5_1, N_67, un1_bckox2_3_net_1, 
        UCK12_RNO_net_1, clk8, clk4, bckox4_sn_N_3, un1_bckox2_1_net_1, 
        bcko;
    
    CFG2 #( .INIT(4'h4) )  master_lrck_inst_1 (.A(cnt_0), .B(i2s_start)
        , .Y(master_lrck));
    CFG4 #( .INIT(16'hF0CA) )  un1_bckox2_3 (.A(clk8), .B(clk4), .C(
        bckox4_sn_N_3), .D(N_68), .Y(un1_bckox2_3_net_1));
    CFG1 #( .INIT(2'h1) )  \cnt_RNO[0]  (.A(\cnt[0]_net_1 ), .Y(
        \cnt_s[0] ));
    SLE \cnt[3]  (.D(\cnt_s[3] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\cnt[3]_net_1 ));
    SLE \cnt[1]  (.D(\cnt_s[1] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\cnt[1]_net_1 ));
    SLE \cnt[5]  (.D(\cnt_s[5]_net_1 ), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(cnt_0));
    CLKINT_PRESERVE UCK10 (.A(bcko), .Y(in_bck_1));
    SLE \cnt[0]  (.D(\cnt_s[0] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\cnt[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  un1_bckox2_1 (.A(bckox2), .B(use_dsd), .Y(
        un1_bckox2_1_net_1));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_s[5]  (.A(VCC_net_1), .B(cnt_0), 
        .C(GND_net_1), .D(GND_net_1), .FCI(\cnt_cry[4]_net_1 ), .S(
        \cnt_s[5]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \cnt_cry[2]  (.A(VCC_net_1), .B(
        \cnt[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_cry[1]_net_1 ), .S(\cnt_s[2] ), .Y(), .FCO(
        \cnt_cry[2]_net_1 ));
    SLE \cnt[4]  (.D(\cnt_s[4] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\cnt[4]_net_1 ));
    SLE \cnt[2]  (.D(\cnt_s[2] ), .CLK(in_bck_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\cnt[2]_net_1 ));
    CFG4 #( .INIT(16'hB931) )  UCK12_RNO (.A(use_dsd), .B(
        un1_bckox2_5_1), .C(N_67), .D(un1_bckox2_3_net_1), .Y(
        UCK12_RNO_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_cry[4]  (.A(VCC_net_1), .B(
        \cnt[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_cry[3]_net_1 ), .S(\cnt_s[4] ), .Y(), .FCO(
        \cnt_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  cnt_s_415 (.A(VCC_net_1), .B(
        \cnt[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(cnt_s_415_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_cry[3]  (.A(VCC_net_1), .B(
        \cnt[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_cry[2]_net_1 ), .S(\cnt_s[3] ), .Y(), .FCO(
        \cnt_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_cry[1]  (.A(VCC_net_1), .B(
        \cnt[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_s_415_FCO), .S(\cnt_s[1] ), .Y(), .FCO(\cnt_cry[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h53) )  UCK12_RNO_0 (.A(N_68), .B(bckox2), .C(
        use_dsd), .Y(un1_bckox2_5_1));
    CLKINT_PRESERVE UCK12 (.A(UCK12_RNO_net_1), .Y(spdif_clock_0));
    CLKINT_PRESERVE UCK14 (.A(un1_bckox2_1_net_1), .Y(dop_clock_0));
    clock_divider UCK0 (.dsd138_ctrl({dsd138_ctrl[2], dsd138_ctrl[1], 
        dsd138_ctrl[0]}), .bcko(bcko), .N_67(N_67), .bckox4_sn_N_3(
        bckox4_sn_N_3), .start_pcm_tx_2(start_pcm_tx_2), .dop_start(
        dop_start), .use_dsd(use_dsd), .i2s_start(i2s_start), .N_68(
        N_68), .bckox2(bckox2), .clk8(clk8), .clk4(clk4), .mclk_1(
        mclk_1), .reset_n_i_i(reset_n_i_i));
    
endmodule


module pcm2dsd(
       dsd138_ctrl,
       cnt_0,
       reset_n_i_i,
       in_bck_1,
       use_dsd,
       i2s_start,
       master_lrck,
       spdif_clock_0,
       dop_clock_0,
       start_pcm_tx_2,
       dop_start,
       mclk_1
    );
input  [2:0] dsd138_ctrl;
output cnt_0;
input  reset_n_i_i;
output in_bck_1;
input  use_dsd;
input  i2s_start;
output master_lrck;
output spdif_clock_0;
output dop_clock_0;
output start_pcm_tx_2;
output dop_start;
input  mclk_1;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    inctrl UIN100 (.dsd138_ctrl({dsd138_ctrl[2], dsd138_ctrl[1], 
        dsd138_ctrl[0]}), .cnt_0(cnt_0), .mclk_1(mclk_1), .dop_start(
        dop_start), .start_pcm_tx_2(start_pcm_tx_2), .dop_clock_0(
        dop_clock_0), .spdif_clock_0(spdif_clock_0), .master_lrck(
        master_lrck), .i2s_start(i2s_start), .use_dsd(use_dsd), 
        .in_bck_1(in_bck_1), .reset_n_i_i(reset_n_i_i));
    GND GND (.Y(GND_net_1));
    
endmodule


module dop_gear(
       dop_right,
       dop_left,
       source_right,
       source_left,
       reset_n_i_3,
       reset_n_i_0_RNIOUJE,
       use_dsd,
       i2s_start,
       reset_n_i_i,
       dop_clock_0
    );
output [15:0] dop_right;
output [15:0] dop_left;
input  [31:0] source_right;
input  [31:0] source_left;
output reset_n_i_3;
input  reset_n_i_0_RNIOUJE;
input  use_dsd;
input  i2s_start;
input  reset_n_i_i;
input  dop_clock_0;

    wire \i[0]_net_1 , VCC_net_1, dop_clock_1, \n_i[0]_net_1 , 
        GND_net_1, \i[1]_net_1 , \i_RNO[1]_net_1 , \i[2]_net_1 , 
        \i_RNO[2]_net_1 , \i[3]_net_1 , \i_RNO[3]_net_1 , 
        \tmp_left[18]_net_1 , n_dop_left_0_sqmuxa_net_1, 
        \tmp_left[19]_net_1 , \tmp_left[20]_net_1 , 
        \tmp_left[21]_net_1 , \tmp_left[22]_net_1 , 
        \tmp_left[23]_net_1 , \tmp_left[24]_net_1 , 
        \tmp_left[25]_net_1 , \tmp_left[26]_net_1 , 
        \tmp_left[27]_net_1 , \tmp_left[28]_net_1 , 
        \tmp_left[29]_net_1 , \tmp_left[30]_net_1 , 
        \tmp_left[31]_net_1 , \tmp_left[3]_net_1 , \tmp_left[4]_net_1 , 
        \tmp_left[5]_net_1 , \tmp_left[6]_net_1 , \tmp_left[7]_net_1 , 
        \tmp_left[8]_net_1 , \tmp_left[9]_net_1 , \tmp_left[10]_net_1 , 
        \tmp_left[11]_net_1 , \tmp_left[12]_net_1 , 
        \tmp_left[13]_net_1 , \tmp_left[14]_net_1 , 
        \tmp_left[15]_net_1 , \tmp_left[16]_net_1 , 
        \tmp_left[17]_net_1 , \tmp_right[20]_net_1 , 
        \tmp_right[21]_net_1 , \tmp_right[22]_net_1 , 
        \tmp_right[23]_net_1 , \tmp_right[24]_net_1 , 
        \tmp_right[25]_net_1 , \tmp_right[26]_net_1 , 
        \tmp_right[27]_net_1 , \tmp_right[28]_net_1 , 
        \tmp_right[29]_net_1 , \tmp_right[30]_net_1 , 
        \tmp_right[31]_net_1 , \tmp_left[0]_net_1 , 
        \tmp_left[1]_net_1 , \tmp_left[2]_net_1 , \tmp_right[5]_net_1 , 
        \tmp_right[6]_net_1 , \tmp_right[7]_net_1 , 
        \tmp_right[8]_net_1 , \tmp_right[9]_net_1 , 
        \tmp_right[10]_net_1 , \tmp_right[11]_net_1 , 
        \tmp_right[12]_net_1 , \tmp_right[13]_net_1 , 
        \tmp_right[14]_net_1 , \tmp_right[15]_net_1 , 
        \tmp_right[16]_net_1 , \tmp_right[17]_net_1 , 
        \tmp_right[18]_net_1 , \tmp_right[19]_net_1 , 
        \n_dop_left[6]_net_1 , n_dop_left_2_sqmuxa_i, 
        \n_dop_left[7]_net_1 , \n_dop_left[8]_net_1 , 
        \n_dop_left[9]_net_1 , \n_dop_left[10]_net_1 , 
        \n_dop_left[11]_net_1 , \n_dop_left[12]_net_1 , 
        \n_dop_left[13]_net_1 , \n_dop_left[14]_net_1 , 
        \n_dop_left[15]_net_1 , \tmp_right[0]_net_1 , 
        \tmp_right[1]_net_1 , \tmp_right[2]_net_1 , 
        \tmp_right[3]_net_1 , \tmp_right[4]_net_1 , 
        \n_dop_right[7]_net_1 , \n_dop_right[8]_net_1 , 
        \n_dop_right[9]_net_1 , \n_dop_right[10]_net_1 , 
        \n_dop_right[11]_net_1 , \n_dop_right[12]_net_1 , 
        \n_dop_right[13]_net_1 , \n_dop_right[14]_net_1 , 
        \n_dop_right[15]_net_1 , \n_dop_left[0]_net_1 , 
        \n_dop_left[1]_net_1 , \n_dop_left[2]_net_1 , 
        \n_dop_left[3]_net_1 , \n_dop_left[4]_net_1 , 
        \n_dop_left[5]_net_1 , \n_dop_right[0]_net_1 , 
        \n_dop_right[1]_net_1 , \n_dop_right[2]_net_1 , 
        \n_dop_right[3]_net_1 , \n_dop_right[4]_net_1 , 
        \n_dop_right[5]_net_1 , \n_dop_right[6]_net_1 , flag_net_1, 
        flag_260_net_1, state_net_1, n_flag6_net_1;
    
    SLE \tmp_left[17]  (.D(source_left[17]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[17]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[12]  (.A(
        \tmp_right[12]_net_1 ), .B(\tmp_right[28]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[12]_net_1 ));
    CFG3 #( .INIT(8'h6A) )  \i_RNO[2]  (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(\i[0]_net_1 ), .Y(\i_RNO[2]_net_1 ));
    SLE \dop_right[6]  (.D(\n_dop_right[6]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[6]));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[6]  (.A(
        \tmp_right[6]_net_1 ), .B(\tmp_right[22]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[6]_net_1 ));
    SLE \tmp_left[26]  (.D(source_left[26]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[26]_net_1 ));
    SLE \tmp_left[13]  (.D(source_left[13]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[13]_net_1 ));
    SLE \tmp_left[1]  (.D(source_left[1]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[1]_net_1 ));
    SLE \tmp_right[15]  (.D(source_right[15]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[15]_net_1 ));
    SLE \tmp_right[7]  (.D(source_right[7]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[7]_net_1 ));
    SLE \dop_left[2]  (.D(\n_dop_left[2]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[2]));
    SLE \tmp_left[14]  (.D(source_left[14]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[14]_net_1 ));
    SLE \tmp_right[29]  (.D(source_right[29]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[29]_net_1 ));
    SLE \i[0]  (.D(\n_i[0]_net_1 ), .CLK(dop_clock_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    SLE \tmp_left[3]  (.D(source_left[3]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[3]_net_1 ));
    CFG4 #( .INIT(16'h6AAA) )  \i_RNO[3]  (.A(\i[3]_net_1 ), .B(
        \i[2]_net_1 ), .C(\i[1]_net_1 ), .D(\i[0]_net_1 ), .Y(
        \i_RNO[3]_net_1 ));
    SLE \tmp_left[5]  (.D(source_left[5]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[5]_net_1 ));
    SLE flag (.D(flag_260_net_1), .CLK(dop_clock_1), .EN(VCC_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(flag_net_1));
    SLE \tmp_left[11]  (.D(source_left[11]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[11]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[11]  (.A(
        \tmp_right[11]_net_1 ), .B(\tmp_right[27]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[11]_net_1 ));
    SLE \dop_right[1]  (.D(\n_dop_right[1]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[1]));
    SLE \dop_right[7]  (.D(\n_dop_right[7]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[7]));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[5]  (.A(\tmp_left[5]_net_1 )
        , .B(\tmp_left[21]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[5]_net_1 ));
    SLE \tmp_right[28]  (.D(source_right[28]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[28]_net_1 ));
    SLE \tmp_left[20]  (.D(source_left[20]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[20]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[8]  (.A(
        \tmp_right[8]_net_1 ), .B(\tmp_right[24]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[8]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[15]  (.A(
        \tmp_right[15]_net_1 ), .B(\tmp_right[31]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[15]_net_1 ));
    SLE \tmp_right[24]  (.D(source_right[24]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[24]_net_1 ));
    SLE \tmp_right[19]  (.D(source_right[19]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[19]_net_1 ));
    CFG2 #( .INIT(4'h8) )  n_dop_left_0_sqmuxa (.A(n_flag6_net_1), .B(
        flag_net_1), .Y(n_dop_left_0_sqmuxa_net_1));
    SLE \dop_left[15]  (.D(\n_dop_left[15]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[15]));
    SLE \dop_right[9]  (.D(\n_dop_right[9]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[9]));
    SLE \dop_right[10]  (.D(\n_dop_right[10]_net_1 ), .CLK(dop_clock_1)
        , .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dop_right[10]));
    SLE \tmp_right[30]  (.D(source_right[30]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[30]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \tmp_left[2]  (.D(source_left[2]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[2]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[14]  (.A(
        \tmp_right[14]_net_1 ), .B(\tmp_right[30]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[14]_net_1 ));
    SLE \dop_right[8]  (.D(\n_dop_right[8]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[8]));
    SLE \dop_right[0]  (.D(\n_dop_right[0]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[0]));
    SLE \tmp_right[18]  (.D(source_right[18]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[18]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[3]  (.A(
        \tmp_right[3]_net_1 ), .B(\tmp_right[19]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[3]_net_1 ));
    SLE \tmp_right[14]  (.D(source_right[14]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[14]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[4]  (.A(
        \tmp_right[4]_net_1 ), .B(\tmp_right[20]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[4]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[9]  (.A(\tmp_left[9]_net_1 )
        , .B(\tmp_left[25]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[9]_net_1 ));
    SLE \tmp_left[22]  (.D(source_left[22]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[22]_net_1 ));
    SLE \tmp_left[27]  (.D(source_left[27]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[27]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \i_RNO[1]  (.A(\i[0]_net_1 ), .B(
        \i[1]_net_1 ), .Y(\i_RNO[1]_net_1 ));
    SLE \dop_left[1]  (.D(\n_dop_left[1]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[1]));
    SLE \tmp_left[23]  (.D(source_left[23]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[23]_net_1 ));
    SLE \dop_left[14]  (.D(\n_dop_left[14]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[14]));
    SLE \tmp_right[2]  (.D(source_right[2]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[2]_net_1 ));
    SLE \dop_left[11]  (.D(\n_dop_left[11]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[11]));
    VCC VCC (.Y(VCC_net_1));
    SLE \tmp_left[24]  (.D(source_left[24]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[24]_net_1 ));
    SLE \tmp_left[18]  (.D(source_left[18]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[18]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[11]  (.A(
        \tmp_left[11]_net_1 ), .B(\tmp_left[27]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_left[11]_net_1 ));
    SLE \tmp_right[26]  (.D(source_right[26]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[26]_net_1 ));
    SLE \dop_left[3]  (.D(\n_dop_left[3]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[3]));
    SLE \dop_left[0]  (.D(\n_dop_left[0]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[0]));
    SLE \tmp_right[31]  (.D(source_right[31]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[31]_net_1 ));
    SLE \tmp_right[5]  (.D(source_right[5]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[5]_net_1 ));
    SLE \tmp_left[8]  (.D(source_left[8]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[8]_net_1 ));
    SLE \tmp_left[21]  (.D(source_left[21]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[21]_net_1 ));
    SLE \tmp_right[9]  (.D(source_right[9]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[9]_net_1 ));
    SLE \dop_left[8]  (.D(\n_dop_left[8]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[8]));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[9]  (.A(
        \tmp_right[9]_net_1 ), .B(\tmp_right[25]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[9]_net_1 ));
    SLE \dop_right[3]  (.D(\n_dop_right[3]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[3]));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[10]  (.A(
        \tmp_left[10]_net_1 ), .B(\tmp_left[26]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_left[10]_net_1 ));
    SLE \tmp_right[3]  (.D(source_right[3]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[3]_net_1 ));
    SLE \tmp_left[19]  (.D(source_left[19]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[19]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[6]  (.A(\tmp_left[6]_net_1 )
        , .B(\tmp_left[22]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[6]_net_1 ));
    SLE \dop_left[4]  (.D(\n_dop_left[4]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[4]));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[5]  (.A(
        \tmp_right[5]_net_1 ), .B(\tmp_right[21]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[5]_net_1 ));
    SLE \tmp_right[16]  (.D(source_right[16]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[16]_net_1 ));
    SLE \tmp_left[9]  (.D(source_left[9]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[9]_net_1 ));
    SLE \dop_right[15]  (.D(\n_dop_right[15]_net_1 ), .CLK(dop_clock_1)
        , .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dop_right[15]));
    SLE \tmp_left[30]  (.D(source_left[30]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[30]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_i[0]  (.A(\i[0]_net_1 ), .B(state_net_1), 
        .Y(\n_i[0]_net_1 ));
    SLE \dop_left[12]  (.D(\n_dop_left[12]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[12]));
    SLE \tmp_right[4]  (.D(source_right[4]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[4]_net_1 ));
    SLE \tmp_right[6]  (.D(source_right[6]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[6]_net_1 ));
    SLE state (.D(VCC_net_1), .CLK(dop_clock_1), .EN(VCC_net_1), .ALn(
        reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(state_net_1));
    SLE \i[2]  (.D(\i_RNO[2]_net_1 ), .CLK(dop_clock_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[0]  (.A(\tmp_left[0]_net_1 )
        , .B(\tmp_left[16]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[0]_net_1 ));
    CLKINT dop_clock_1_RNO (.A(dop_clock_0), .Y(dop_clock_1));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[12]  (.A(
        \tmp_left[12]_net_1 ), .B(\tmp_left[28]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_left[12]_net_1 ));
    SLE \dop_left[5]  (.D(\n_dop_left[5]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[5]));
    SLE \tmp_right[22]  (.D(source_right[22]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[22]_net_1 ));
    SLE \dop_right[11]  (.D(\n_dop_right[11]_net_1 ), .CLK(dop_clock_1)
        , .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dop_right[11]));
    SLE \dop_right[14]  (.D(\n_dop_right[14]_net_1 ), .CLK(dop_clock_1)
        , .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dop_right[14]));
    SLE \tmp_left[28]  (.D(source_left[28]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[28]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[13]  (.A(
        \tmp_left[13]_net_1 ), .B(\tmp_left[29]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_left[13]_net_1 ));
    SLE \tmp_right[20]  (.D(source_right[20]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[20]_net_1 ));
    CFG3 #( .INIT(8'h08) )  reset_n_i (.A(i2s_start), .B(use_dsd), .C(
        reset_n_i_0_RNIOUJE), .Y(reset_n_i_3));
    SLE \tmp_right[27]  (.D(source_right[27]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[27]_net_1 ));
    SLE \tmp_left[6]  (.D(source_left[6]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[6]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[7]  (.A(\tmp_left[7]_net_1 )
        , .B(\tmp_left[23]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[7]_net_1 ));
    SLE \dop_left[6]  (.D(\n_dop_left[6]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[6]));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[13]  (.A(
        \tmp_right[13]_net_1 ), .B(\tmp_right[29]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[13]_net_1 ));
    SLE \tmp_left[15]  (.D(source_left[15]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[15]_net_1 ));
    SLE \tmp_left[29]  (.D(source_left[29]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[29]_net_1 ));
    SLE \tmp_right[12]  (.D(source_right[12]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[12]_net_1 ));
    SLE \dop_right[5]  (.D(\n_dop_right[5]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[5]));
    SLE \tmp_right[10]  (.D(source_right[10]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[10]_net_1 ));
    SLE \tmp_right[8]  (.D(source_right[8]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[8]_net_1 ));
    SLE \tmp_left[16]  (.D(source_left[16]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[16]_net_1 ));
    SLE \dop_right[13]  (.D(\n_dop_right[13]_net_1 ), .CLK(dop_clock_1)
        , .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dop_right[13]));
    SLE \tmp_right[17]  (.D(source_right[17]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[17]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[8]  (.A(\tmp_left[8]_net_1 )
        , .B(\tmp_left[24]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[8]_net_1 ));
    SLE \dop_left[10]  (.D(\n_dop_left[10]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[10]));
    SLE \tmp_left[31]  (.D(source_left[31]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[31]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[10]  (.A(
        \tmp_right[10]_net_1 ), .B(\tmp_right[26]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[10]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[4]  (.A(\tmp_left[4]_net_1 )
        , .B(\tmp_left[20]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[4]_net_1 ));
    SLE \tmp_right[23]  (.D(source_right[23]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[23]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  n_flag6 (.A(\i[3]_net_1 ), .B(
        \i[2]_net_1 ), .C(\i[1]_net_1 ), .D(\i[0]_net_1 ), .Y(
        n_flag6_net_1));
    SLE \tmp_right[1]  (.D(source_right[1]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[1]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[3]  (.A(\tmp_left[3]_net_1 )
        , .B(\tmp_left[19]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[3]_net_1 ));
    SLE \dop_right[4]  (.D(\n_dop_right[4]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[4]));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[14]  (.A(
        \tmp_left[14]_net_1 ), .B(\tmp_left[30]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_left[14]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_left[2]  (.A(\tmp_left[2]_net_1 )
        , .B(\tmp_left[18]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[2]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[0]  (.A(
        \tmp_right[0]_net_1 ), .B(\tmp_right[16]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[0]_net_1 ));
    SLE \dop_right[12]  (.D(\n_dop_right[12]_net_1 ), .CLK(dop_clock_1)
        , .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dop_right[12]));
    SLE \tmp_right[21]  (.D(source_right[21]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[21]_net_1 ));
    SLE \tmp_left[4]  (.D(source_left[4]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[4]_net_1 ));
    SLE \tmp_left[10]  (.D(source_left[10]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[10]_net_1 ));
    CFG2 #( .INIT(4'hB) )  state_RNIC1DQ (.A(n_flag6_net_1), .B(
        state_net_1), .Y(n_dop_left_2_sqmuxa_i));
    SLE \tmp_right[13]  (.D(source_right[13]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[13]_net_1 ));
    SLE \tmp_left[7]  (.D(source_left[7]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[7]_net_1 ));
    SLE \i[3]  (.D(\i_RNO[3]_net_1 ), .CLK(dop_clock_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    CFG4 #( .INIT(16'hAFCF) )  \n_dop_right[2]  (.A(
        \tmp_right[2]_net_1 ), .B(\tmp_right[18]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[2]_net_1 ));
    SLE \dop_left[7]  (.D(\n_dop_left[7]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[7]));
    SLE \tmp_right[0]  (.D(source_right[0]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[0]_net_1 ));
    SLE \dop_right[2]  (.D(\n_dop_right[2]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_right[2]));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[15]  (.A(
        \tmp_left[15]_net_1 ), .B(\tmp_left[31]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_left[15]_net_1 ));
    SLE \i[1]  (.D(\i_RNO[1]_net_1 ), .CLK(dop_clock_1), .EN(VCC_net_1)
        , .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG3 #( .INIT(8'h4A) )  flag_260 (.A(n_flag6_net_1), .B(
        state_net_1), .C(flag_net_1), .Y(flag_260_net_1));
    SLE \dop_left[13]  (.D(\n_dop_left[13]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[13]));
    SLE \tmp_right[11]  (.D(source_right[11]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[11]_net_1 ));
    SLE \dop_left[9]  (.D(\n_dop_left[9]_net_1 ), .CLK(dop_clock_1), 
        .EN(n_dop_left_2_sqmuxa_i), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dop_left[9]));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[1]  (.A(
        \tmp_right[1]_net_1 ), .B(\tmp_right[17]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[1]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_left[1]  (.A(\tmp_left[1]_net_1 )
        , .B(\tmp_left[17]_net_1 ), .C(n_flag6_net_1), .D(flag_net_1), 
        .Y(\n_dop_left[1]_net_1 ));
    SLE \tmp_right[25]  (.D(source_right[25]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_right[25]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \n_dop_right[7]  (.A(
        \tmp_right[7]_net_1 ), .B(\tmp_right[23]_net_1 ), .C(
        n_flag6_net_1), .D(flag_net_1), .Y(\n_dop_right[7]_net_1 ));
    SLE \tmp_left[12]  (.D(source_left[12]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[12]_net_1 ));
    SLE \tmp_left[0]  (.D(source_left[0]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[0]_net_1 ));
    SLE \tmp_left[25]  (.D(source_left[25]), .CLK(dop_clock_1), .EN(
        n_dop_left_0_sqmuxa_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tmp_left[25]_net_1 ));
    
endmodule


module crc16(
       crc0,
       bits_0,
       crc_en,
       sdclk_n_1,
       crc_clr_i
    );
output [14:0] crc0;
input  bits_0;
input  crc_en;
input  sdclk_n_1;
input  crc_clr_i;

    wire VCC_net_1, GND_net_1, N_62_i, \CRC[15]_net_1 , inv, N_63_i;
    
    SLE \CRC[10]  (.D(crc0[9]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[10]));
    SLE \CRC[0]  (.D(inv), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[0]));
    SLE \CRC[2]  (.D(crc0[1]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[2]));
    SLE \CRC[14]  (.D(crc0[13]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[14]));
    SLE \CRC[13]  (.D(crc0[12]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[13]));
    GND GND (.Y(GND_net_1));
    SLE \CRC[5]  (.D(N_63_i), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[5]));
    CFG2 #( .INIT(4'h6) )  inv_i_o3 (.A(bits_0), .B(\CRC[15]_net_1 ), 
        .Y(inv));
    CFG2 #( .INIT(4'h6) )  \CRCX_1_i_0_x2[12]  (.A(inv), .B(crc0[11]), 
        .Y(N_62_i));
    SLE \CRC[1]  (.D(crc0[0]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[1]));
    SLE \CRC[6]  (.D(crc0[5]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[6]));
    SLE \CRC[7]  (.D(crc0[6]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[7]));
    SLE \CRC[3]  (.D(crc0[2]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[3]));
    SLE \CRC[12]  (.D(N_62_i), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[12]));
    CFG2 #( .INIT(4'h6) )  \CRCX_1_0_a3_0_x2[5]  (.A(inv), .B(crc0[4]), 
        .Y(N_63_i));
    SLE \CRC[9]  (.D(crc0[8]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[9]));
    SLE \CRC[11]  (.D(crc0[10]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[11]));
    SLE \CRC[4]  (.D(crc0[3]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[4]));
    SLE \CRC[15]  (.D(crc0[14]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\CRC[15]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \CRC[8]  (.D(crc0[7]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc0[8]));
    
endmodule


module crc16_0(
       crc1,
       bits_0,
       crc_en,
       sdclk_n_1,
       crc_clr_i
    );
output [14:0] crc1;
input  bits_0;
input  crc_en;
input  sdclk_n_1;
input  crc_clr_i;

    wire VCC_net_1, GND_net_1, \CRCX_1[12] , \CRC[15]_net_1 , inv, 
        \CRCX_1[5] ;
    
    SLE \CRC[10]  (.D(crc1[9]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[10]));
    SLE \CRC[0]  (.D(inv), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[0]));
    SLE \CRC[2]  (.D(crc1[1]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[2]));
    SLE \CRC[14]  (.D(crc1[13]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[14]));
    SLE \CRC[13]  (.D(crc1[12]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[13]));
    GND GND (.Y(GND_net_1));
    SLE \CRC[5]  (.D(\CRCX_1[5] ), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[5]));
    CFG3 #( .INIT(8'h96) )  \CRCX_1_i[12]  (.A(bits_0), .B(crc1[11]), 
        .C(\CRC[15]_net_1 ), .Y(\CRCX_1[12] ));
    CFG2 #( .INIT(4'h6) )  inv_i_o3 (.A(bits_0), .B(\CRC[15]_net_1 ), 
        .Y(inv));
    SLE \CRC[1]  (.D(crc1[0]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[1]));
    SLE \CRC[6]  (.D(crc1[5]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[6]));
    SLE \CRC[7]  (.D(crc1[6]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[7]));
    SLE \CRC[3]  (.D(crc1[2]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[3]));
    SLE \CRC[12]  (.D(\CRCX_1[12] ), .CLK(sdclk_n_1), .EN(crc_en), 
        .ALn(crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(crc1[12]));
    SLE \CRC[9]  (.D(crc1[8]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[9]));
    CFG3 #( .INIT(8'h96) )  \CRCX_1_0_a3[5]  (.A(bits_0), .B(crc1[4]), 
        .C(\CRC[15]_net_1 ), .Y(\CRCX_1[5] ));
    SLE \CRC[11]  (.D(crc1[10]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[11]));
    SLE \CRC[4]  (.D(crc1[3]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[4]));
    SLE \CRC[15]  (.D(crc1[14]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\CRC[15]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \CRC[8]  (.D(crc1[7]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc1[8]));
    
endmodule


module crc16_1(
       crc2,
       bits_0,
       crc_en,
       sdclk_n_1,
       crc_clr_i
    );
output [14:0] crc2;
input  bits_0;
input  crc_en;
input  sdclk_n_1;
input  crc_clr_i;

    wire VCC_net_1, GND_net_1, \CRCX_1[12] , \CRC[15]_net_1 , inv, 
        \CRCX_1[5] ;
    
    SLE \CRC[10]  (.D(crc2[9]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[10]));
    SLE \CRC[0]  (.D(inv), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[0]));
    SLE \CRC[2]  (.D(crc2[1]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[2]));
    SLE \CRC[14]  (.D(crc2[13]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[14]));
    SLE \CRC[13]  (.D(crc2[12]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[13]));
    GND GND (.Y(GND_net_1));
    SLE \CRC[5]  (.D(\CRCX_1[5] ), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[5]));
    CFG3 #( .INIT(8'h96) )  \CRCX_1_i[12]  (.A(bits_0), .B(crc2[11]), 
        .C(\CRC[15]_net_1 ), .Y(\CRCX_1[12] ));
    CFG2 #( .INIT(4'h6) )  inv_i_o3 (.A(bits_0), .B(\CRC[15]_net_1 ), 
        .Y(inv));
    SLE \CRC[1]  (.D(crc2[0]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[1]));
    SLE \CRC[6]  (.D(crc2[5]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[6]));
    SLE \CRC[7]  (.D(crc2[6]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[7]));
    SLE \CRC[3]  (.D(crc2[2]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[3]));
    SLE \CRC[12]  (.D(\CRCX_1[12] ), .CLK(sdclk_n_1), .EN(crc_en), 
        .ALn(crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(crc2[12]));
    SLE \CRC[9]  (.D(crc2[8]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[9]));
    CFG3 #( .INIT(8'h96) )  \CRCX_1_0_a3[5]  (.A(bits_0), .B(crc2[4]), 
        .C(\CRC[15]_net_1 ), .Y(\CRCX_1[5] ));
    SLE \CRC[11]  (.D(crc2[10]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[11]));
    SLE \CRC[4]  (.D(crc2[3]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[4]));
    SLE \CRC[15]  (.D(crc2[14]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\CRC[15]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \CRC[8]  (.D(crc2[7]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc2[8]));
    
endmodule


module crc16_2(
       crc3,
       bits_0,
       crc_en,
       sdclk_n_1,
       crc_clr_i
    );
output [14:0] crc3;
input  bits_0;
input  crc_en;
input  sdclk_n_1;
input  crc_clr_i;

    wire VCC_net_1, GND_net_1, N_82_i, \CRC[15]_net_1 , inv, N_83_i;
    
    SLE \CRC[10]  (.D(crc3[9]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[10]));
    CFG3 #( .INIT(8'h96) )  \CRCX_1_0_a3_0_x4[5]  (.A(bits_0), .B(
        crc3[4]), .C(\CRC[15]_net_1 ), .Y(N_83_i));
    SLE \CRC[0]  (.D(inv), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[0]));
    SLE \CRC[2]  (.D(crc3[1]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[2]));
    SLE \CRC[14]  (.D(crc3[13]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[14]));
    SLE \CRC[13]  (.D(crc3[12]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[13]));
    GND GND (.Y(GND_net_1));
    SLE \CRC[5]  (.D(N_83_i), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[5]));
    CFG2 #( .INIT(4'h6) )  inv_i_o3 (.A(bits_0), .B(\CRC[15]_net_1 ), 
        .Y(inv));
    SLE \CRC[1]  (.D(crc3[0]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[1]));
    SLE \CRC[6]  (.D(crc3[5]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[6]));
    SLE \CRC[7]  (.D(crc3[6]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[7]));
    SLE \CRC[3]  (.D(crc3[2]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[3]));
    SLE \CRC[12]  (.D(N_82_i), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[12]));
    SLE \CRC[9]  (.D(crc3[8]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[9]));
    SLE \CRC[11]  (.D(crc3[10]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[11]));
    SLE \CRC[4]  (.D(crc3[3]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[4]));
    SLE \CRC[15]  (.D(crc3[14]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\CRC[15]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \CRCX_1_i_0_x4[12]  (.A(bits_0), .B(
        crc3[11]), .C(\CRC[15]_net_1 ), .Y(N_82_i));
    SLE \CRC[8]  (.D(crc3[7]), .CLK(sdclk_n_1), .EN(crc_en), .ALn(
        crc_clr_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(crc3[8]));
    
endmodule


module sd_data(
       total_blocks,
       sd_data_out,
       din,
       sd_data_in,
       status_0,
       in_cmd,
       sd_read_start,
       sd_write_start,
       data_bus_busy,
       wen,
       is_last_data,
       sdclk_n_1,
       sdclk_n_i,
       u8_sb_0_HPMS_READY,
       data_out_en_ret_fast_i,
       sd_data_out_en_i_i
    );
input  [3:0] total_blocks;
output [3:0] sd_data_out;
output [31:0] din;
input  [3:0] sd_data_in;
input  status_0;
input  in_cmd;
input  sd_read_start;
input  sd_write_start;
output data_bus_busy;
output wen;
output is_last_data;
input  sdclk_n_1;
input  sdclk_n_i;
input  u8_sb_0_HPMS_READY;
output data_out_en_ret_fast_i;
output sd_data_out_en_i_i;

    wire crc_clr_net_1, crc_clr_0, sd_data_out_en_i, 
        data_out_en_ret_fast_net_1, crc_clr_i, \data0[3]_net_1 , 
        VCC_net_1, GND_net_1, \odin[22]_net_1 , N_64_i, N_388_i, 
        \odin[23]_net_1 , N_3458_i, \odin[24]_net_1 , N_3457_i, 
        \odin[25]_net_1 , N_3456_i, \odin[26]_net_1 , N_3455_i, 
        \odin[27]_net_1 , \n_din[27]_net_1 , \blkn[0]_net_1 , 
        \n_blkn[0]_net_1 , \blkn[1]_net_1 , \n_blkn[1]_net_1 , 
        \blkn[2]_net_1 , N_3770_i, \blkn[3]_net_1 , N_3769_i, 
        \data0[0]_net_1 , \data0[1]_net_1 , \data0[2]_net_1 , 
        \odin[7]_net_1 , N_68_i, \odin[8]_net_1 , N_66_i, 
        \odin[9]_net_1 , \n_din[9] , \odin[10]_net_1 , 
        \n_din[10]_net_1 , \odin[11]_net_1 , \n_din[11]_net_1 , 
        \odin[12]_net_1 , \n_din[12] , \odin[13]_net_1 , 
        \n_din[13]_net_1 , \odin[14]_net_1 , \n_din[14]_net_1 , 
        \odin[15]_net_1 , \n_din[15]_net_1 , \odin[16]_net_1 , 
        \n_din[16] , \odin[17]_net_1 , \n_din[17] , \odin[18]_net_1 , 
        \n_din[18]_net_1 , \odin[19]_net_1 , \n_din[19]_net_1 , 
        \odin[20]_net_1 , \n_din[20]_net_1 , \odin[21]_net_1 , 
        \n_din[21] , \n_AX[28] , un1_n_data_bus_busy8_2_i, \n_AX[29] , 
        \n_AX[30] , \n_AX[31] , \dq[0]_net_1 , dq_148_net_1, 
        \dq[1]_net_1 , dq_149_net_1, \dq[2]_net_1 , dq_150_net_1, 
        \dq[3]_net_1 , dq_151_net_1, \odin[0]_net_1 , \n_din[0] , 
        \odin[1]_net_1 , \n_din[1] , \odin[2]_net_1 , N_72_i, 
        \odin[3]_net_1 , \n_din[3]_net_1 , \odin[4]_net_1 , \n_din[4] , 
        \odin[5]_net_1 , \n_din[5] , \odin[6]_net_1 , N_70_i, 
        \n_AX[13] , \n_AX[14] , \n_AX[15] , \n_AX[16] , \n_AX[17] , 
        \n_AX[18] , \n_AX[19] , \n_AX[20] , \n_AX[21] , \n_AX[22] , 
        \n_AX[23] , \n_AX[24] , \n_AX[25] , \n_AX[26] , \n_AX[27] , 
        \bits[2]_net_1 , \bits_ldmx[2]_net_1 , 
        n_data_out_en_3_sqmuxa_i, \bits[3]_net_1 , 
        \bits_ldmx[3]_net_1 , N_3767_i, N_3768_i, \n_AX[2] , \n_AX[3] , 
        \n_AX[4] , \n_AX[5] , \n_AX[6] , \n_AX[7] , \n_AX[8] , 
        \n_AX[9] , \n_AX[10] , \n_AX[11] , \n_AX[12] , 
        \n_data_out_iv_i_0[0]_net_1 , un1_state_9_i, 
        \n_data_out_iv_i_0[1]_net_1 , \n_data_out_iv_i_0[2]_net_1 , 
        \n_data_out_iv_i_0[3]_net_1 , \bits[0]_net_1 , 
        \bits_ldmx_4_1_0_wmux_0_Y[0] , \bits[1]_net_1 , 
        \bits_ldmx[1]_net_1 , n_crc_clr_iv_i, un1_state_19_i, 
        n_is_last_data_iv_i, N_384_i, n_AX_0_sqmuxa_net_1, N_387_i, 
        N_383_i, crc_en_net_1, \state[6]_net_1 , N_379_i, 
        \state[5]_net_1 , \state_ns[5] , N_692_i, \state[7]_net_1 , 
        \state_ns[7] , \state[0]_net_1 , \state_ns[0] , 
        \state[1]_net_1 , \state_ns[1] , \state[2]_net_1 , N_687_i, 
        \state[3]_net_1 , \state_ns[3] , \state[4]_net_1 , 
        \state_ns[4] , \i[0]_net_1 , \i_lm[0] , N_3446_i, \i[1]_net_1 , 
        \i_lm[1] , \i[2]_net_1 , \i_lm[2] , \i[3]_net_1 , \i_lm[3] , 
        \i[4]_net_1 , \i_lm[4] , \i[5]_net_1 , \i_lm[5] , \i[6]_net_1 , 
        \i_lm[6] , \i[7]_net_1 , \i_lm[7] , \i[8]_net_1 , \i_lm[8] , 
        \i[9]_net_1 , \i_lm[9] , sd_data_out_eni, un1_state_6_i, 
        i_s_417_FCO, \i_cry[1]_net_1 , \i_s[1] , \i_cry[2]_net_1 , 
        \i_s[2] , \i_cry[3]_net_1 , \i_s[3] , \i_cry[4]_net_1 , 
        \i_s[4] , \i_cry[5]_net_1 , \i_s[5] , \i_cry[6]_net_1 , 
        \i_s[6] , \i_cry[7]_net_1 , \i_s[7] , \i_s[9]_net_1 , 
        \i_cry[8]_net_1 , \i_s[8] , \bits_en[0]_net_1 , 
        \bits_ldmx_2[0]_net_1 , N_3934_i, \bits_ldmx_4_1_0_y0[0] , 
        \bits_ldmx_4_1_0_co0[0] , \bits_ldmx_0[0]_net_1 , 
        n_bits_sn_N_11_mux, N_793, \crc3[5] , \crc3[4] , 
        \n_bits_10_0_0_y0[3] , \n_bits_10_0_0_co0[3] , \crc3[13] , 
        \crc3[12] , N_800, \crc2[8] , \crc2[0] , \n_bits_12_0_0_y0[2] , 
        \n_bits_12_0_0_co0[2] , \crc2[9] , \crc2[1] , N_792, \crc2[5] , 
        \crc2[4] , \n_bits_10_0_0_y0[2] , \n_bits_10_0_0_co0[2] , 
        \crc2[13] , \crc2[12] , N_801, \crc3[8] , \crc3[0] , 
        \n_bits_12_0_0_y0[3] , \n_bits_12_0_0_co0[3] , \crc3[9] , 
        \crc3[1] , N_3947, \crc1[5] , \crc1[4] , 
        \n_bits_10_i_m2_0_0_y0[1] , \n_bits_10_i_m2_0_0_co0[1] , 
        \crc1[13] , \crc1[12] , N_3780, \crc1[6] , \crc1[2] , 
        \n_bits_13_i_m3_0_0_y0[1] , \n_bits_13_i_m3_0_0_co0[1] , 
        \crc1[7] , \crc1[3] , N_3779, \crc2[6] , \crc2[2] , 
        \n_bits_13_i_m3_0_0_y0[2] , \n_bits_13_i_m3_0_0_co0[2] , 
        \crc2[7] , \crc2[3] , N_3946, \crc0[8] , \crc0[0] , 
        \n_bits_12_i_m2_0_0_y0[0] , \n_bits_12_i_m2_0_0_co0[0] , 
        \crc0[9] , \crc0[1] , N_3945, \crc1[8] , \crc1[0] , 
        \n_bits_12_i_m2_0_0_y0[1] , \n_bits_12_i_m2_0_0_co0[1] , 
        \crc1[9] , \crc1[1] , N_3944, \crc0[6] , \crc0[2] , 
        \n_bits_13_i_m2_0_0_y0[0] , \n_bits_13_i_m2_0_0_co0[0] , 
        \crc0[7] , \crc0[3] , N_3778, \crc3[6] , \crc3[2] , 
        \n_bits_13_i_m3_0_0_y0[3] , \n_bits_13_i_m3_0_0_co0[3] , 
        \crc3[7] , \crc3[3] , un48_n_i_c4, n_i_sn_N_8_mux, 
        \n_i_0_iv_0_1[4]_net_1 , \state_ns_0_a2_0_RNI7N2R[5]_net_1 , 
        un1_state_21_i, \i_lm_0_1_0[0]_net_1 , n_i_iv_0_a2_out, 
        \n_i_iv_0_a2_2_0[0]_net_1 , n_i_sn_N_7_mux, N_789, 
        \bits_ldmx_1[3]_net_1 , N_818, N_788, \bits_ldmx_1[2]_net_1 , 
        N_817, N_787, \bits_ldmx_1[1]_net_1 , N_816, CO2_1, CO2, 
        \n_i_0_iv_0[4]_net_1 , \crc1[10] , \n_bits_11_i_m3_1[1]_net_1 , 
        N_3782, \crc1[11] , \crc1[14] , \crc0[12] , 
        \n_bits_16_i_m2_1_1[0]_net_1 , N_3941, \crc0[13] , \crc0[14] , 
        \crc2[10] , \n_bits_11_i_m3_1[2]_net_1 , N_3781, \crc2[11] , 
        \crc2[14] , \crc3[10] , \n_bits_15_i_m4_1[3]_net_1 , N_3791, 
        \crc3[11] , \crc3[14] , \n_bits_16_bm[3]_net_1 , 
        \n_bits_16_am[3]_net_1 , \n_bits_16_bm[2]_net_1 , 
        \n_bits_16_am[2]_net_1 , \n_bits_16_bm[1]_net_1 , 
        \n_bits_16_am[1]_net_1 , n_bits_17_sqmuxa, \n_dq_0[3]_net_1 , 
        \n_dq_0[0]_net_1 , \n_dq_0[1]_net_1 , \n_dq_0[2]_net_1 , 
        \state_ns_0_o4_1[3]_net_1 , un1_i_4lt4, 
        un1_state_16_i_a2_0_net_1, n_i_0_iv_0_a2_0_out_0, 
        n_i_0_iv_0_a2_0_out, un48_n_i_axbxc1_net_1, 
        n_data_out_1_sqmuxa_1_net_1, N_3935_i, N_4074, N_3968_1, 
        n_wen7_net_1, N_702_i, N_78, N_137, N_386_i, \crc0[10] , 
        \crc0[11] , N_3937, \crc0[4] , \crc0[5] , N_3936, 
        un1_state_18_1_net_1, n_is_last_data6_4_net_1, 
        n_is_last_data6_3_0_net_1, \state_ns_0_a2_0_1_1_a2_1[5]_net_1 , 
        N_700, n_data_out6_net_1, n_dq8, N_3819, N_378, N_3971, 
        un48_n_i_axbxc2_net_1, un1_state_21_0_0_1_net_1, 
        \n_bits_16_i_1[0]_net_1 , n_data_out_2_sqmuxa_1_net_1, N_3970, 
        N_702, un48_n_i_axbxc3_net_1, N_135, N_726, N_719, N_76_i, 
        n_i_0_iv_0_a2_out, \state_ns_0_0[0]_net_1 , 
        \state_ns_0_0[1]_net_1 , un1_state_21_0_0_2_net_1, 
        \n_bits_16_i_0[0]_net_1 , n_data_out_2_sqmuxa_2_net_1, N_729, 
        N_731, n_is_last_data6_net_1, un1_n_blkn_0_sqmuxa_net_1, 
        \state_ns_i_0[6]_net_1 , \n_i_0_iv_0_a2_0[2]_net_1 , 
        \n_i_0_iv_0_a2_0[3]_net_1 , n_i_0_iv_0_a2_1_out, CO1, 
        \n_i_0_iv_0[1]_net_1 , un1_state_21_0_0_5_net_1, 
        \n_i_0_iv_0[5]_net_1 ;
    
    SLE \odin[2]  (.D(N_72_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[2]_net_1 ));
    SLE \AX[30]  (.D(\n_AX[30] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[30]));
    SLE \state[0]  (.D(\state_ns[0] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_10_0_0_wmux_0[3]  (.A(
        \n_bits_10_0_0_y0[3] ), .B(\i[3]_net_1 ), .C(\crc3[5] ), .D(
        \crc3[4] ), .FCI(\n_bits_10_0_0_co0[3] ), .S(), .Y(N_793), 
        .FCO());
    CFG4 #( .INIT(16'hA060) )  \n_i_0_iv_0_a2_s[1]  (.A(\i[1]_net_1 ), 
        .B(\i[0]_net_1 ), .C(\state[4]_net_1 ), .D(status_0), .Y(
        n_i_0_iv_0_a2_out));
    SLE \odin[8]  (.D(N_66_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[8]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \n_bits_16_am[1]  (.A(\i[3]_net_1 ), .B(
        N_3782), .C(N_3780), .Y(\n_bits_16_am[1]_net_1 ));
    CFG3 #( .INIT(8'h53) )  \n_bits_11_i_m3_1[2]  (.A(\crc2[11] ), .B(
        \crc2[14] ), .C(\i[2]_net_1 ), .Y(\n_bits_11_i_m3_1[2]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \n_bits_16_ns[2]  (.A(\i[1]_net_1 ), .B(
        \n_bits_16_bm[2]_net_1 ), .C(\n_bits_16_am[2]_net_1 ), .Y(
        N_817));
    SLE \i[7]  (.D(\i_lm[7] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_13_i_m3_0_0_wmux[1]  (.A(
        \i[2]_net_1 ), .B(\i[0]_net_1 ), .C(\crc1[7] ), .D(\crc1[3] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_13_i_m3_0_0_y0[1] ), .FCO(
        \n_bits_13_i_m3_0_0_co0[1] ));
    CFG3 #( .INIT(8'h53) )  \n_bits_11_i_m3_1[1]  (.A(\crc1[11] ), .B(
        \crc1[14] ), .C(\i[2]_net_1 ), .Y(\n_bits_11_i_m3_1[1]_net_1 ));
    SLE \blkn[2]  (.D(N_3770_i), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\blkn[2]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \bits_ldmx_4_1_0_wmux[0]  (.A(
        n_bits_sn_N_11_mux), .B(\bits_en[0]_net_1 ), .C(
        \bits_ldmx_0[0]_net_1 ), .D(\bits[0]_net_1 ), .FCI(VCC_net_1), 
        .S(), .Y(\bits_ldmx_4_1_0_y0[0] ), .FCO(
        \bits_ldmx_4_1_0_co0[0] ));
    SLE \AX[10]  (.D(\n_AX[10] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[10]));
    CFG3 #( .INIT(8'hB8) )  \n_bits_9[2]  (.A(din[30]), .B(
        \state[6]_net_1 ), .C(n_bits_17_sqmuxa), .Y(N_788));
    CFG1 #( .INIT(2'h1) )  data_out_en_ret_fast_RNI3LM5 (.A(
        data_out_en_ret_fast_net_1), .Y(data_out_en_ret_fast_i));
    CFG2 #( .INIT(4'h8) )  \n_i_0_iv_0_a2_0_s[3]  (.A(\i[3]_net_1 ), 
        .B(\state[4]_net_1 ), .Y(n_i_0_iv_0_a2_0_out_0));
    SLE \i[0]  (.D(\i_lm[0] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_13_i_m3_0_0_wmux_0[2]  (.A(
        \n_bits_13_i_m3_0_0_y0[2] ), .B(\i[0]_net_1 ), .C(\crc2[6] ), 
        .D(\crc2[2] ), .FCI(\n_bits_13_i_m3_0_0_co0[2] ), .S(), .Y(
        N_3779), .FCO());
    SLE \state[6]  (.D(N_692_i), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[6]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[9]  (.A(\state[0]_net_1 ), .B(
        \odin[5]_net_1 ), .Y(\n_din[9] ));
    SLE \AX[17]  (.D(\n_AX[17] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[17]));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[25]  (.A(\state[0]_net_1 ), .B(
        \odin[21]_net_1 ), .Y(N_3456_i));
    CFG2 #( .INIT(4'h4) )  \n_din[10]  (.A(\state[0]_net_1 ), .B(
        \odin[6]_net_1 ), .Y(\n_din[10]_net_1 ));
    CFG4 #( .INIT(16'hCECA) )  \n_i_0_iv_0_a2_0[2]  (.A(
        n_i_0_iv_0_a2_0_out), .B(un48_n_i_axbxc2_net_1), .C(
        n_i_sn_N_7_mux), .D(\n_i_iv_0_a2_2_0[0]_net_1 ), .Y(
        \n_i_0_iv_0_a2_0[2]_net_1 ));
    SLE \data0[3]  (.D(sd_data_in[3]), .CLK(sdclk_n_i), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\data0[3]_net_1 ));
    CFG4 #( .INIT(16'hCBC8) )  \bits_ldmx_2[0]  (.A(din[28]), .B(
        \state[6]_net_1 ), .C(n_bits_sn_N_11_mux), .D(n_bits_17_sqmuxa)
        , .Y(\bits_ldmx_2[0]_net_1 ));
    SLE \AX[20]  (.D(\n_AX[20] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[20]));
    CFG4 #( .INIT(16'hD888) )  \i_lm_0[2]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(\i_s[2] ), .C(
        un1_state_21_i), .D(\n_i_0_iv_0_a2_0[2]_net_1 ), .Y(\i_lm[2] ));
    CFG4 #( .INIT(16'hFFEF) )  \state_ns_0_o4[3]  (.A(\i[0]_net_1 ), 
        .B(\state_ns_0_o4_1[3]_net_1 ), .C(\i[4]_net_1 ), .D(
        \i[3]_net_1 ), .Y(N_702));
    CFG4 #( .INIT(16'h006C) )  \blkn_RNO[3]  (.A(\blkn[2]_net_1 ), .B(
        \blkn[3]_net_1 ), .C(CO1), .D(\state[0]_net_1 ), .Y(N_3769_i));
    CFG4 #( .INIT(16'hEEF0) )  dq_149 (.A(\n_dq_0[1]_net_1 ), .B(
        N_3819), .C(\dq[1]_net_1 ), .D(N_378), .Y(dq_149_net_1));
    SLE \AX[4]  (.D(\n_AX[4] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[4]));
    CFG2 #( .INIT(4'h8) )  un1_n_data_out_1_sqmuxa_RNO (.A(status_0), 
        .B(\state[4]_net_1 ), .Y(N_3935_i));
    crc16 UCRC0 (.crc0({\crc0[14] , \crc0[13] , \crc0[12] , \crc0[11] , 
        \crc0[10] , \crc0[9] , \crc0[8] , \crc0[7] , \crc0[6] , 
        \crc0[5] , \crc0[4] , \crc0[3] , \crc0[2] , \crc0[1] , 
        \crc0[0] }), .bits_0(\bits[0]_net_1 ), .crc_en(crc_en_net_1), 
        .sdclk_n_1(sdclk_n_1), .crc_clr_i(crc_clr_i));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_13_i_m2_0_0_wmux[0]  (.A(
        \i[2]_net_1 ), .B(\i[0]_net_1 ), .C(\crc0[7] ), .D(\crc0[3] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_13_i_m2_0_0_y0[0] ), .FCO(
        \n_bits_13_i_m2_0_0_co0[0] ));
    SLE \odin[7]  (.D(N_68_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[7]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \n_bits_16_bm[3]  (.A(N_801), .B(
        \i[2]_net_1 ), .C(N_793), .Y(\n_bits_16_bm[3]_net_1 ));
    SLE \AX[27]  (.D(\n_AX[27] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[27]));
    crc16_0 UCRC1 (.crc1({\crc1[14] , \crc1[13] , \crc1[12] , 
        \crc1[11] , \crc1[10] , \crc1[9] , \crc1[8] , \crc1[7] , 
        \crc1[6] , \crc1[5] , \crc1[4] , \crc1[3] , \crc1[2] , 
        \crc1[1] , \crc1[0] }), .bits_0(\bits[1]_net_1 ), .crc_en(
        crc_en_net_1), .sdclk_n_1(sdclk_n_1), .crc_clr_i(crc_clr_i));
    SLE \data_out[1]  (.D(\n_data_out_iv_i_0[1]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_9_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sd_data_out[1]));
    CFG3 #( .INIT(8'hB8) )  \n_bits_16_i_m2_0[0]  (.A(\crc0[10] ), .B(
        \i[0]_net_1 ), .C(\crc0[11] ), .Y(N_3937));
    CFG4 #( .INIT(16'hFFFE) )  un1_state_21_0_0_5 (.A(n_i_sn_N_8_mux), 
        .B(n_i_sn_N_7_mux), .C(un1_state_21_0_0_2_net_1), .D(N_729), 
        .Y(un1_state_21_0_0_5_net_1));
    CFG4 #( .INIT(16'h80BF) )  \n_bits_11_i_m3[1]  (.A(\crc1[10] ), .B(
        \i[2]_net_1 ), .C(\i[0]_net_1 ), .D(
        \n_bits_11_i_m3_1[1]_net_1 ), .Y(N_3782));
    CFG4 #( .INIT(16'h0001) )  \bits_en[0]  (.A(\state[4]_net_1 ), .B(
        \state[0]_net_1 ), .C(N_729), .D(N_378), .Y(\bits_en[0]_net_1 )
        );
    SLE \AX[12]  (.D(\n_AX[12] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[12]));
    CFG4 #( .INIT(16'hCCEA) )  \n_i_0_iv_0[1]  (.A(n_i_0_iv_0_a2_out), 
        .B(un48_n_i_axbxc1_net_1), .C(\n_i_iv_0_a2_2_0[0]_net_1 ), .D(
        n_i_sn_N_7_mux), .Y(\n_i_0_iv_0[1]_net_1 ));
    CFG4 #( .INIT(16'h0A0B) )  \n_data_out_iv_i_0[2]  (.A(
        \bits[2]_net_1 ), .B(\state[6]_net_1 ), .C(N_4074), .D(
        n_i_sn_N_8_mux), .Y(\n_data_out_iv_i_0[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  un48_n_i_axbxc1 (.A(\i[0]_net_1 ), .B(
        \i[1]_net_1 ), .Y(un48_n_i_axbxc1_net_1));
    SLE \state[4]  (.D(\state_ns[4] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[4]_net_1 ));
    CFG2 #( .INIT(4'hD) )  crc_en_RNO (.A(un1_state_16_i_a2_0_net_1), 
        .B(\state[6]_net_1 ), .Y(N_379_i));
    CFG4 #( .INIT(16'h0010) )  \state_ns_0_o4_1_RNIBD8Q[3]  (.A(
        \i[0]_net_1 ), .B(\state_ns_0_o4_1[3]_net_1 ), .C(\i[4]_net_1 )
        , .D(\i[3]_net_1 ), .Y(N_702_i));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[2]  (.A(\state[0]_net_1 ), .B(
        \dq[2]_net_1 ), .Y(N_72_i));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h4) )  \n_din[27]  (.A(\state[0]_net_1 ), .B(
        \odin[23]_net_1 ), .Y(\n_din[27]_net_1 ));
    SLE \state[7]  (.D(\state_ns[7] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[7]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_12_0_0_wmux[3]  (.A(
        \i[3]_net_1 ), .B(\i[0]_net_1 ), .C(\crc3[9] ), .D(\crc3[1] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_12_0_0_y0[3] ), .FCO(
        \n_bits_12_0_0_co0[3] ));
    CFG3 #( .INIT(8'hD8) )  \n_bits_16_ns[3]  (.A(\i[1]_net_1 ), .B(
        \n_bits_16_bm[3]_net_1 ), .C(\n_bits_16_am[3]_net_1 ), .Y(
        N_818));
    SLE \dq[3]  (.D(dq_151_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\dq[3]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \n_bits_16_am[3]  (.A(\i[3]_net_1 ), .B(
        N_3791), .C(N_3778), .Y(\n_bits_16_am[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  data_out_en_ret_RNIMJB9 (.A(
        sd_data_out_en_i), .Y(sd_data_out_en_i_i));
    SLE \state[5]  (.D(\state_ns[5] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[5]_net_1 ));
    SLE \AX[22]  (.D(\n_AX[22] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[22]));
    CFG2 #( .INIT(4'h8) )  n_AX_0_sqmuxa (.A(n_wen7_net_1), .B(
        \state[2]_net_1 ), .Y(n_AX_0_sqmuxa_net_1));
    CFG2 #( .INIT(4'h4) )  \n_din[3]  (.A(\state[0]_net_1 ), .B(
        \dq[3]_net_1 ), .Y(\n_din[3]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_13_i_m3_0_0_wmux[3]  (.A(
        \i[2]_net_1 ), .B(\i[0]_net_1 ), .C(\crc3[7] ), .D(\crc3[3] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_13_i_m3_0_0_y0[3] ), .FCO(
        \n_bits_13_i_m3_0_0_co0[3] ));
    CFG4 #( .INIT(16'h3A33) )  \bits_ldmx[3]  (.A(N_789), .B(
        \bits_ldmx_1[3]_net_1 ), .C(n_bits_sn_N_11_mux), .D(
        \bits_en[0]_net_1 ), .Y(\bits_ldmx[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \state_ns_i_o2[6]  (.A(\state[6]_net_1 ), 
        .B(n_is_last_data6_net_1), .C(n_i_sn_N_8_mux), .Y(
        \state_ns[7] ));
    SLE \AX[13]  (.D(\n_AX[13] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[13]));
    CFG4 #( .INIT(16'hFEF0) )  un1_state_21_0_0_2 (.A(\dq[0]_net_1 ), 
        .B(\dq[1]_net_1 ), .C(un1_state_21_0_0_1_net_1), .D(
        \state[1]_net_1 ), .Y(un1_state_21_0_0_2_net_1));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[4]  (.A(din[0]), .B(
        \odin[0]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(\n_AX[4] )
        );
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[6]  (.A(din[2]), .B(
        \odin[2]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(\n_AX[6] )
        );
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[1]  (.A(\state[0]_net_1 ), .B(
        \dq[1]_net_1 ), .Y(\n_din[1] ));
    CFG2 #( .INIT(4'hB) )  n_AX_1_sqmuxa_1_i_o2 (.A(n_wen7_net_1), .B(
        \state[6]_net_1 ), .Y(N_78));
    CFG3 #( .INIT(8'hB8) )  \n_bits_16_bm[2]  (.A(N_800), .B(
        \i[2]_net_1 ), .C(N_792), .Y(\n_bits_16_bm[2]_net_1 ));
    SLE \odin[20]  (.D(\n_din[20]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[20]_net_1 ));
    SLE \dq[2]  (.D(dq_150_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\dq[2]_net_1 ));
    SLE \odin[10]  (.D(\n_din[10]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[10]_net_1 ));
    SLE \AX[14]  (.D(\n_AX[14] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[14]));
    SLE \data_out[2]  (.D(\n_data_out_iv_i_0[2]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_9_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sd_data_out[2]));
    CFG3 #( .INIT(8'hFE) )  \state_RNIR6VD[3]  (.A(\state[3]_net_1 ), 
        .B(\state[2]_net_1 ), .C(\state[0]_net_1 ), .Y(N_384_i));
    CFG4 #( .INIT(16'h0002) )  n_data_out6 (.A(\i[4]_net_1 ), .B(
        \i[3]_net_1 ), .C(\i[2]_net_1 ), .D(\i[0]_net_1 ), .Y(
        n_data_out6_net_1));
    CFG3 #( .INIT(8'hB8) )  \n_bits_9[3]  (.A(din[31]), .B(
        \state[6]_net_1 ), .C(n_bits_17_sqmuxa), .Y(N_789));
    CFG2 #( .INIT(4'h4) )  \n_din[13]  (.A(\state[0]_net_1 ), .B(
        \odin[9]_net_1 ), .Y(\n_din[13]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_10_0_0_wmux_0[2]  (.A(
        \n_bits_10_0_0_y0[2] ), .B(\i[3]_net_1 ), .C(\crc2[5] ), .D(
        \crc2[4] ), .FCI(\n_bits_10_0_0_co0[2] ), .S(), .Y(N_792), 
        .FCO());
    SLE \AX[23]  (.D(\n_AX[23] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[23]));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[12]  (.A(\state[0]_net_1 ), .B(
        \odin[8]_net_1 ), .Y(\n_din[12] ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[19]  (.A(din[15]), .B(
        \odin[15]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[19] ));
    SLE \dq[1]  (.D(dq_149_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\dq[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \state_RNI0HTU[3]  (.A(N_702_i), .B(
        \state[3]_net_1 ), .Y(n_i_sn_N_7_mux));
    CFG4 #( .INIT(16'h0008) )  \n_bits_16_i_a2_1[0]  (.A(\i[3]_net_1 ), 
        .B(\i[1]_net_1 ), .C(N_3936), .D(\i[2]_net_1 ), .Y(N_3970));
    SLE \bits[1]  (.D(\bits_ldmx[1]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_data_out_en_3_sqmuxa_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\bits[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \bits_ldmx_0[0]  (.A(n_bits_sn_N_11_mux), 
        .B(\bits[0]_net_1 ), .C(\state[6]_net_1 ), .Y(
        \bits_ldmx_0[0]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[26]  (.A(din[22]), .B(
        \odin[22]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[26] ));
    CFG4 #( .INIT(16'hFF04) )  \n_bits_16_i_1[0]  (.A(\i[1]_net_1 ), 
        .B(\i[3]_net_1 ), .C(N_3944), .D(N_3971), .Y(
        \n_bits_16_i_1[0]_net_1 ));
    SLE \AX[31]  (.D(\n_AX[31] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[31]));
    CFG3 #( .INIT(8'h08) )  n_data_out_2_sqmuxa_2 (.A(
        n_data_out_2_sqmuxa_1_net_1), .B(\state[3]_net_1 ), .C(
        n_data_out6_net_1), .Y(n_data_out_2_sqmuxa_2_net_1));
    SLE \i[9]  (.D(\i_lm[9] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    SLE \AX[24]  (.D(\n_AX[24] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[24]));
    CFG4 #( .INIT(16'hCE0A) )  un1_n_blkn_0_sqmuxa (.A(
        \state[1]_net_1 ), .B(\state[6]_net_1 ), .C(N_700), .D(
        n_is_last_data6_net_1), .Y(un1_n_blkn_0_sqmuxa_net_1));
    CFG2 #( .INIT(4'h8) )  \n_i_0_iv_0_a2_0_s[2]  (.A(\i[2]_net_1 ), 
        .B(\state[4]_net_1 ), .Y(n_i_0_iv_0_a2_0_out));
    CFG3 #( .INIT(8'hE4) )  \n_bits_16_am[2]  (.A(\i[3]_net_1 ), .B(
        N_3781), .C(N_3779), .Y(\n_bits_16_am[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \AX_RNO[1]  (.A(\state[2]_net_1 ), .B(
        \dq[1]_net_1 ), .Y(N_3768_i));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[25]  (.A(din[21]), .B(
        \odin[21]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[25] ));
    CFG2 #( .INIT(4'h8) )  \AX_RNO[2]  (.A(\state[2]_net_1 ), .B(
        \dq[2]_net_1 ), .Y(\n_AX[2] ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hE) )  un1_n_data_out_1_sqmuxa (.A(
        n_data_out_1_sqmuxa_1_net_1), .B(N_3935_i), .Y(N_4074));
    CFG4 #( .INIT(16'hDDDC) )  un1_state_21_0_0 (.A(
        n_is_last_data6_net_1), .B(un1_state_21_0_0_5_net_1), .C(
        \state[2]_net_1 ), .D(\state[6]_net_1 ), .Y(un1_state_21_i));
    CFG4 #( .INIT(16'hECA0) )  \state_ns_0[3]  (.A(\state[2]_net_1 ), 
        .B(\state[3]_net_1 ), .C(n_is_last_data6_net_1), .D(N_702), .Y(
        \state_ns[3] ));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[8]  (.A(\state[0]_net_1 ), .B(
        \odin[4]_net_1 ), .Y(N_66_i));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_12_0_0_wmux_0[3]  (.A(
        \n_bits_12_0_0_y0[3] ), .B(\i[0]_net_1 ), .C(\crc3[8] ), .D(
        \crc3[0] ), .FCI(\n_bits_12_0_0_co0[3] ), .S(), .Y(N_801), 
        .FCO());
    CFG4 #( .INIT(16'h3A33) )  \bits_ldmx[1]  (.A(N_787), .B(
        \bits_ldmx_1[1]_net_1 ), .C(n_bits_sn_N_11_mux), .D(
        \bits_en[0]_net_1 ), .Y(\bits_ldmx[1]_net_1 ));
    SLE \AX[11]  (.D(\n_AX[11] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[11]));
    CFG4 #( .INIT(16'hF4F0) )  \state_ns_0[5]  (.A(sd_write_start), .B(
        sd_read_start), .C(N_729), .D(\state[0]_net_1 ), .Y(
        \state_ns[5] ));
    CFG2 #( .INIT(4'h1) )  \n_bits_16_i_a2_0_2[0]  (.A(\i[2]_net_1 ), 
        .B(\i[3]_net_1 ), .Y(un1_i_4lt4));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[22]  (.A(\state[0]_net_1 ), .B(
        \odin[18]_net_1 ), .Y(N_64_i));
    CFG4 #( .INIT(16'hF1F0) )  \state_ns_0_0[0]  (.A(sd_write_start), 
        .B(sd_read_start), .C(N_719), .D(\state[0]_net_1 ), .Y(
        \state_ns_0_0[0]_net_1 ));
    SLE \odin[24]  (.D(N_3457_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[24]_net_1 ));
    CFG4 #( .INIT(16'hEEF0) )  dq_150 (.A(\n_dq_0[2]_net_1 ), .B(
        N_3819), .C(\dq[2]_net_1 ), .D(N_378), .Y(dq_150_net_1));
    SLE \data0[1]  (.D(sd_data_in[1]), .CLK(sdclk_n_i), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\data0[1]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \n_dq_0[0]  (.A(\data0[0]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\n_dq_0[0]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[9]  (.A(din[5]), .B(
        \odin[5]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(\n_AX[9] )
        );
    SLE \odin[14]  (.D(\n_din[14]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[14]_net_1 ));
    SLE \odin[26]  (.D(N_3455_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[26]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \n_blkn[1]  (.A(\blkn[0]_net_1 ), .B(
        \blkn[1]_net_1 ), .C(un1_n_blkn_0_sqmuxa_net_1), .D(
        \state[0]_net_1 ), .Y(\n_blkn[1]_net_1 ));
    CFG3 #( .INIT(8'h0D) )  \n_bits_16_i_a2_0_2_RNIDD0G[0]  (.A(
        \i[4]_net_1 ), .B(un1_i_4lt4), .C(\i[5]_net_1 ), .Y(N_135));
    SLE \odin[16]  (.D(\n_din[16] ), .CLK(sdclk_n_1), .EN(N_388_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\odin[16]_net_1 ));
    SLE crc_clr (.D(n_crc_clr_iv_i), .CLK(sdclk_n_1), .EN(
        un1_state_19_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(crc_clr_0)
        );
    SLE \odin[27]  (.D(\n_din[27]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[27]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[23]  (.A(din[19]), .B(
        \odin[19]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[23] ));
    SLE \odin[17]  (.D(\n_din[17] ), .CLK(sdclk_n_1), .EN(N_388_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\odin[17]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \n_bits_16_ns[1]  (.A(\i[1]_net_1 ), .B(
        \n_bits_16_bm[1]_net_1 ), .C(\n_bits_16_am[1]_net_1 ), .Y(
        N_816));
    SLE \odin[18]  (.D(\n_din[18]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[18]_net_1 ));
    SLE \AX[21]  (.D(\n_AX[21] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[21]));
    SLE \odin[25]  (.D(N_3456_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[25]_net_1 ));
    CFG4 #( .INIT(16'h0A4E) )  \state_RNO[2]  (.A(\state[1]_net_1 ), 
        .B(\state[2]_net_1 ), .C(N_700), .D(n_is_last_data6_net_1), .Y(
        N_687_i));
    CFG4 #( .INIT(16'h0A0B) )  \n_data_out_iv_i_0[3]  (.A(
        \bits[3]_net_1 ), .B(\state[6]_net_1 ), .C(N_4074), .D(
        n_i_sn_N_8_mux), .Y(\n_data_out_iv_i_0[3]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[27]  (.A(din[23]), .B(
        \odin[23]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[27] ));
    CLKINT crc_clr_RNI1MED (.A(crc_clr_0), .Y(crc_clr_net_1));
    CFG4 #( .INIT(16'h0A8E) )  \n_dq8_1.CO2_1  (.A(total_blocks[1]), 
        .B(total_blocks[0]), .C(\blkn[1]_net_1 ), .D(\blkn[0]_net_1 ), 
        .Y(CO2_1));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[28]  (.A(din[24]), .B(
        \odin[24]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[28] ));
    SLE \odin[15]  (.D(\n_din[15]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[15]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \AX_RNO[3]  (.A(\state[2]_net_1 ), .B(
        \dq[3]_net_1 ), .Y(\n_AX[3] ));
    SLE \AX[3]  (.D(\n_AX[3] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[3]));
    SLE \blkn[0]  (.D(\n_blkn[0]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \blkn[0]_net_1 ));
    SLE \AX[9]  (.D(\n_AX[9] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[9]));
    CFG4 #( .INIT(16'h6AAA) )  un48_n_i_axbxc3 (.A(\i[3]_net_1 ), .B(
        \i[1]_net_1 ), .C(\i[0]_net_1 ), .D(\i[2]_net_1 ), .Y(
        un48_n_i_axbxc3_net_1));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[23]  (.A(\state[0]_net_1 ), .B(
        \odin[19]_net_1 ), .Y(N_3458_i));
    CFG3 #( .INIT(8'h4C) )  crc_clr_RNO (.A(N_76_i), .B(N_386_i), .C(
        n_dq8), .Y(n_crc_clr_iv_i));
    CFG4 #( .INIT(16'h000D) )  \state_RNO[6]  (.A(\state[7]_net_1 ), 
        .B(n_dq8), .C(\state_ns_i_0[6]_net_1 ), .D(\state_ns[7] ), .Y(
        N_692_i));
    CFG3 #( .INIT(8'hAC) )  \n_bits_16_i_m2[0]  (.A(\crc0[4] ), .B(
        \crc0[5] ), .C(\i[0]_net_1 ), .Y(N_3936));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[0]  (.A(\state[0]_net_1 ), .B(
        \dq[0]_net_1 ), .Y(\n_din[0] ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_12_i_m2_0_0_wmux[0]  (.A(
        \i[3]_net_1 ), .B(\i[0]_net_1 ), .C(\crc0[9] ), .D(\crc0[1] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_12_i_m2_0_0_y0[0] ), .FCO(
        \n_bits_12_i_m2_0_0_co0[0] ));
    CFG4 #( .INIT(16'hD888) )  \i_lm_0[3]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(\i_s[3] ), .C(
        un1_state_21_i), .D(\n_i_0_iv_0_a2_0[3]_net_1 ), .Y(\i_lm[3] ));
    SLE wen_inst_1 (.D(n_AX_0_sqmuxa_net_1), .CLK(sdclk_n_1), .EN(
        N_384_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(wen));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_10_0_0_wmux[2]  (.A(
        \i[0]_net_1 ), .B(\i[3]_net_1 ), .C(\crc2[13] ), .D(\crc2[12] )
        , .FCI(VCC_net_1), .S(), .Y(\n_bits_10_0_0_y0[2] ), .FCO(
        \n_bits_10_0_0_co0[2] ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[5]  (.A(din[1]), .B(
        \odin[1]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(\n_AX[5] )
        );
    CFG4 #( .INIT(16'h0D00) )  \n_bits_16_i_a2_0_2_RNI6LLK[0]  (.A(
        \i[4]_net_1 ), .B(un1_i_4lt4), .C(\i[5]_net_1 ), .D(
        \state[7]_net_1 ), .Y(n_i_sn_N_8_mux));
    CFG4 #( .INIT(16'hEEF0) )  dq_151 (.A(\n_dq_0[3]_net_1 ), .B(
        N_3819), .C(\dq[3]_net_1 ), .D(N_378), .Y(dq_151_net_1));
    SLE \odin[21]  (.D(\n_din[21] ), .CLK(sdclk_n_1), .EN(N_388_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\odin[21]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[18]  (.A(din[14]), .B(
        \odin[14]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[18] ));
    SLE \odin[11]  (.D(\n_din[11]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[11]_net_1 ));
    SLE \odin[23]  (.D(N_3458_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[23]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \n_dq_0[3]  (.A(\data0[3]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\n_dq_0[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[6]_net_1 ), .S(\i_s[7] ), .Y(), .FCO(\i_cry[7]_net_1 ));
    CFG4 #( .INIT(16'h0015) )  crc_clr_RNO_0 (.A(n_bits_sn_N_11_mux), 
        .B(un1_state_16_i_a2_0_net_1), .C(N_386_i), .D(N_729), .Y(
        un1_state_19_i));
    crc16_1 UCRC2 (.crc2({\crc2[14] , \crc2[13] , \crc2[12] , 
        \crc2[11] , \crc2[10] , \crc2[9] , \crc2[8] , \crc2[7] , 
        \crc2[6] , \crc2[5] , \crc2[4] , \crc2[3] , \crc2[2] , 
        \crc2[1] , \crc2[0] }), .bits_0(\bits[2]_net_1 ), .crc_en(
        crc_en_net_1), .sdclk_n_1(sdclk_n_1), .crc_clr_i(crc_clr_i));
    CFG3 #( .INIT(8'h20) )  \n_bits_16_i_a2_2[0]  (.A(\i[2]_net_1 ), 
        .B(N_3946), .C(\i[1]_net_1 ), .Y(N_3971));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[15]  (.A(din[11]), .B(
        \odin[11]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[15] ));
    SLE \odin[0]  (.D(\n_din[0] ), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[0]_net_1 ));
    CFG3 #( .INIT(8'h8E) )  \n_dq8_1.CO3  (.A(CO2), .B(total_blocks[3])
        , .C(\blkn[3]_net_1 ), .Y(n_dq8));
    SLE \odin[13]  (.D(\n_din[13]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[13]_net_1 ));
    CFG3 #( .INIT(8'hFB) )  \state_RNIQ37I2[7]  (.A(n_dq8), .B(
        \state[7]_net_1 ), .C(N_135), .Y(n_data_out_en_3_sqmuxa_i));
    CFG4 #( .INIT(16'h2000) )  \state_ns_i_a2_0[6]  (.A(N_137), .B(
        \state[6]_net_1 ), .C(un1_i_4lt4), .D(
        \state_ns_0_a2_0_1_1_a2_1[5]_net_1 ), .Y(N_731));
    CFG4 #( .INIT(16'hEA40) )  \i_lm_0[6]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(un1_state_21_i), .C(
        \i[6]_net_1 ), .D(\i_s[6] ), .Y(\i_lm[6] ));
    CFG4 #( .INIT(16'hEEF0) )  dq_148 (.A(\n_dq_0[0]_net_1 ), .B(
        N_3819), .C(\dq[0]_net_1 ), .D(N_378), .Y(dq_148_net_1));
    SLE data_out_en_ret_fast (.D(sd_data_out_eni), .CLK(sdclk_n_1), 
        .EN(un1_state_6_i), .ALn(u8_sb_0_HPMS_READY), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        data_out_en_ret_fast_net_1));
    CFG4 #( .INIT(16'h8000) )  un48_n_i_ac0_5 (.A(\i[3]_net_1 ), .B(
        \i[1]_net_1 ), .C(\i[0]_net_1 ), .D(\i[2]_net_1 ), .Y(
        un48_n_i_c4));
    CFG4 #( .INIT(16'hCECA) )  \n_i_0_iv_0_a2_0[3]  (.A(
        n_i_0_iv_0_a2_0_out_0), .B(un48_n_i_axbxc3_net_1), .C(
        n_i_sn_N_7_mux), .D(\n_i_iv_0_a2_2_0[0]_net_1 ), .Y(
        \n_i_0_iv_0_a2_0[3]_net_1 ));
    SLE \i[2]  (.D(\i_lm[2] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    CFG4 #( .INIT(16'h0A0B) )  \n_data_out_iv_i_0[1]  (.A(
        \bits[1]_net_1 ), .B(\state[6]_net_1 ), .C(N_4074), .D(
        n_i_sn_N_8_mux), .Y(\n_data_out_iv_i_0[1]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \n_dq_0[1]  (.A(\data0[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\n_dq_0[1]_net_1 ));
    SLE \blkn[3]  (.D(N_3769_i), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\blkn[3]_net_1 ));
    CFG4 #( .INIT(16'hF0F2) )  \n_bits_16_i_0[0]  (.A(N_3968_1), .B(
        \i[1]_net_1 ), .C(N_3970), .D(N_3937), .Y(
        \n_bits_16_i_0[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \state_ns_i_a4_0_a2[6]  (.A(
        \state[7]_net_1 ), .B(\i[4]_net_1 ), .C(\i[5]_net_1 ), .Y(
        n_bits_sn_N_11_mux));
    CFG3 #( .INIT(8'h53) )  \n_bits_15_i_m4_1[3]  (.A(\crc3[11] ), .B(
        \crc3[14] ), .C(\i[2]_net_1 ), .Y(\n_bits_15_i_m4_1[3]_net_1 ));
    SLE \odin[19]  (.D(\n_din[19]_net_1 ), .CLK(sdclk_n_1), .EN(
        N_388_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \odin[19]_net_1 ));
    SLE \dq[0]  (.D(dq_148_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\dq[0]_net_1 ));
    SLE crc_en (.D(\state[6]_net_1 ), .CLK(sdclk_n_1), .EN(N_379_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(crc_en_net_1));
    CFG4 #( .INIT(16'h153F) )  \state_ns_0_o4_RNIP8GV[1]  (.A(
        \state[1]_net_1 ), .B(in_cmd), .C(N_729), .D(N_700), .Y(
        N_3446_i));
    CFG4 #( .INIT(16'h0040) )  \state_ns_0_a2_2[0]  (.A(\i[1]_net_1 ), 
        .B(\i[0]_net_1 ), .C(\state[4]_net_1 ), .D(status_0), .Y(N_719)
        );
    CFG4 #( .INIT(16'hD888) )  \i_lm_0[1]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(\i_s[1] ), .C(
        un1_state_21_i), .D(\n_i_0_iv_0[1]_net_1 ), .Y(\i_lm[1] ));
    CFG3 #( .INIT(8'h53) )  \bits_ldmx_1[2]  (.A(N_817), .B(
        \bits[2]_net_1 ), .C(\bits_en[0]_net_1 ), .Y(
        \bits_ldmx_1[2]_net_1 ));
    SLE \AX[0]  (.D(N_3767_i), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[0]));
    CFG4 #( .INIT(16'h0001) )  \state_ns_0_a2_0_1_1_a2_1[5]  (.A(
        \i[7]_net_1 ), .B(\i[6]_net_1 ), .C(\i[5]_net_1 ), .D(
        \i[4]_net_1 ), .Y(\state_ns_0_a2_0_1_1_a2_1[5]_net_1 ));
    SLE data_out_en_ret (.D(sd_data_out_eni), .CLK(sdclk_n_1), .EN(
        un1_state_6_i), .ALn(u8_sb_0_HPMS_READY), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sd_data_out_en_i));
    SLE \data_out[3]  (.D(\n_data_out_iv_i_0[3]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_9_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sd_data_out[3]));
    CFG2 #( .INIT(4'h1) )  un1_state_16_i_a2_0 (.A(\state[0]_net_1 ), 
        .B(\state[7]_net_1 ), .Y(un1_state_16_i_a2_0_net_1));
    CFG4 #( .INIT(16'hF0FE) )  \state_ns_0_a2_0_RNI7N2R[5]  (.A(
        \state[6]_net_1 ), .B(\state[2]_net_1 ), .C(N_729), .D(
        n_is_last_data6_net_1), .Y(\state_ns_0_a2_0_RNI7N2R[5]_net_1 ));
    CFG4 #( .INIT(16'h333B) )  un1_state_18 (.A(\state[7]_net_1 ), .B(
        un1_state_18_1_net_1), .C(N_135), .D(n_dq8), .Y(
        sd_data_out_eni));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[24]  (.A(\state[0]_net_1 ), .B(
        \odin[20]_net_1 ), .Y(N_3457_i));
    CFG2 #( .INIT(4'h4) )  \n_din[14]  (.A(\state[0]_net_1 ), .B(
        \odin[10]_net_1 ), .Y(\n_din[14]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[22]  (.A(din[18]), .B(
        \odin[18]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[22] ));
    CFG4 #( .INIT(16'h3F5F) )  n_data_out_2_sqmuxa_1 (.A(N_3968_1), .B(
        un1_i_4lt4), .C(\i[4]_net_1 ), .D(\i[1]_net_1 ), .Y(
        n_data_out_2_sqmuxa_1_net_1));
    SLE \state[3]  (.D(\state_ns[3] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[3]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[16]  (.A(din[12]), .B(
        \odin[12]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[16] ));
    SLE \bits[2]  (.D(\bits_ldmx[2]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_data_out_en_3_sqmuxa_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\bits[2]_net_1 ));
    CFG4 #( .INIT(16'hF0B0) )  \state_ns_0_a2[4]  (.A(\i[1]_net_1 ), 
        .B(\i[0]_net_1 ), .C(\state[4]_net_1 ), .D(status_0), .Y(N_726)
        );
    CFG4 #( .INIT(16'h0AB2) )  \n_i_0_iv_0_1[4]  (.A(un48_n_i_c4), .B(
        n_i_sn_N_8_mux), .C(\i[4]_net_1 ), .D(\state[4]_net_1 ), .Y(
        \n_i_0_iv_0_1[4]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[11]  (.A(din[7]), .B(
        \odin[7]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[11] ));
    CFG4 #( .INIT(16'h80BF) )  \n_bits_11_i_m3[2]  (.A(\crc2[10] ), .B(
        \i[2]_net_1 ), .C(\i[0]_net_1 ), .D(
        \n_bits_11_i_m3_1[2]_net_1 ), .Y(N_3781));
    SLE \AX[19]  (.D(\n_AX[19] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[19]));
    CFG4 #( .INIT(16'h8000) )  n_is_last_data6_4 (.A(\i[4]_net_1 ), .B(
        \i[5]_net_1 ), .C(\i[3]_net_1 ), .D(\i[1]_net_1 ), .Y(
        n_is_last_data6_4_net_1));
    SLE \AX[15]  (.D(\n_AX[15] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[15]));
    SLE \odin[1]  (.D(\n_din[1] ), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[1]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_12_i_m2_0_0_wmux_0[0]  (.A(
        \n_bits_12_i_m2_0_0_y0[0] ), .B(\i[0]_net_1 ), .C(\crc0[8] ), 
        .D(\crc0[0] ), .FCI(\n_bits_12_i_m2_0_0_co0[0] ), .S(), .Y(
        N_3946), .FCO());
    CFG1 #( .INIT(2'h1) )  crc_clr_RNI1MED_0 (.A(crc_clr_net_1), .Y(
        crc_clr_i));
    SLE \AX[18]  (.D(\n_AX[18] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[18]));
    SLE \i[6]  (.D(\i_lm[6] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    CFG4 #( .INIT(16'h3A33) )  \bits_ldmx[2]  (.A(N_788), .B(
        \bits_ldmx_1[2]_net_1 ), .C(n_bits_sn_N_11_mux), .D(
        \bits_en[0]_net_1 ), .Y(\bits_ldmx[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(i_s_417_FCO), 
        .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    CFG4 #( .INIT(16'hAAAE) )  \state_ns_0[4]  (.A(N_726), .B(
        \state[3]_net_1 ), .C(n_dq8), .D(N_702), .Y(\state_ns[4] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[4]  (.D(\i_lm[4] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    SLE \odin[9]  (.D(\n_din[9] ), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[9]_net_1 ));
    CFG2 #( .INIT(4'h8) )  n_bits_17_sqmuxa_0_a2 (.A(n_i_sn_N_8_mux), 
        .B(\i[4]_net_1 ), .Y(n_bits_17_sqmuxa));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(\i_cry[6]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \state_RNI63A9[2]  (.A(\state[0]_net_1 ), 
        .B(\state[2]_net_1 ), .Y(N_388_i));
    CFG3 #( .INIT(8'h47) )  \n_bits_16_i_m2_1_1[0]  (.A(\crc0[13] ), 
        .B(\i[1]_net_1 ), .C(\crc0[14] ), .Y(
        \n_bits_16_i_m2_1_1[0]_net_1 ));
    SLE data_bus_busy_inst_1 (.D(N_387_i), .CLK(sdclk_n_1), .EN(
        N_383_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(data_bus_busy));
    CFG4 #( .INIT(16'hCCCE) )  \state_ns_0[0]  (.A(\state[7]_net_1 ), 
        .B(\state_ns_0_0[0]_net_1 ), .C(N_135), .D(n_dq8), .Y(
        \state_ns[0] ));
    SLE \odin[3]  (.D(\n_din[3]_net_1 ), .CLK(sdclk_n_1), .EN(N_388_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\odin[3]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[17]  (.A(din[13]), .B(
        \odin[13]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[17] ));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[26]  (.A(\state[0]_net_1 ), .B(
        \odin[22]_net_1 ), .Y(N_3455_i));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_13_i_m3_0_0_wmux[2]  (.A(
        \i[2]_net_1 ), .B(\i[0]_net_1 ), .C(\crc2[7] ), .D(\crc2[3] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_13_i_m3_0_0_y0[2] ), .FCO(
        \n_bits_13_i_m3_0_0_co0[2] ));
    CFG4 #( .INIT(16'hEA40) )  \i_lm_0[8]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(un1_state_21_i), .C(
        \i[8]_net_1 ), .D(\i_s[8] ), .Y(\i_lm[8] ));
    SLE \AX[29]  (.D(\n_AX[29] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[29]));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_12_0_0_wmux_0[2]  (.A(
        \n_bits_12_0_0_y0[2] ), .B(\i[0]_net_1 ), .C(\crc2[8] ), .D(
        \crc2[0] ), .FCI(\n_bits_12_0_0_co0[2] ), .S(), .Y(N_800), 
        .FCO());
    SLE \AX[25]  (.D(\n_AX[25] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[25]));
    SLE \AX[28]  (.D(\n_AX[28] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[28]));
    CFG2 #( .INIT(4'h4) )  \n_din[18]  (.A(\state[0]_net_1 ), .B(
        \odin[14]_net_1 ), .Y(\n_din[18]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \n_i_iv_0_a2_2_0[0]  (.A(n_i_sn_N_8_mux), 
        .B(\state[4]_net_1 ), .Y(\n_i_iv_0_a2_2_0[0]_net_1 ));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_12_i_m2_0_0_wmux_0[1]  (.A(
        \n_bits_12_i_m2_0_0_y0[1] ), .B(\i[0]_net_1 ), .C(\crc1[8] ), 
        .D(\crc1[0] ), .FCI(\n_bits_12_i_m2_0_0_co0[1] ), .S(), .Y(
        N_3945), .FCO());
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[7]  (.A(din[3]), .B(
        \odin[3]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(\n_AX[7] )
        );
    CFG4 #( .INIT(16'h8000) )  n_is_last_data6_3_0 (.A(\i[9]_net_1 ), 
        .B(\i[8]_net_1 ), .C(\i[7]_net_1 ), .D(\i[6]_net_1 ), .Y(
        n_is_last_data6_3_0_net_1));
    SLE \AX[6]  (.D(\n_AX[6] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[6]));
    CFG3 #( .INIT(8'h6A) )  un48_n_i_axbxc2 (.A(\i[2]_net_1 ), .B(
        \i[0]_net_1 ), .C(\i[1]_net_1 ), .Y(un48_n_i_axbxc2_net_1));
    CFG4 #( .INIT(16'h0A0B) )  \n_data_out_iv_i_0[0]  (.A(
        \bits[0]_net_1 ), .B(\state[6]_net_1 ), .C(N_4074), .D(
        n_i_sn_N_8_mux), .Y(\n_data_out_iv_i_0[0]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \n_bits_16_i_a2_0_1[0]  (.A(\i[2]_net_1 ), 
        .B(\i[3]_net_1 ), .Y(N_3968_1));
    SLE \bits[0]  (.D(\bits_ldmx_4_1_0_wmux_0_Y[0] ), .CLK(sdclk_n_1), 
        .EN(n_data_out_en_3_sqmuxa_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\bits[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \AX_RNO[0]  (.A(\state[2]_net_1 ), .B(
        \dq[0]_net_1 ), .Y(N_3767_i));
    CFG2 #( .INIT(4'h1) )  \state_ns_i_a2_1_0[6]  (.A(\state[6]_net_1 )
        , .B(\state[5]_net_1 ), .Y(N_386_i));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[14]  (.A(din[10]), .B(
        \odin[10]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[14] ));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[5]  (.A(\state[0]_net_1 ), .B(
        \odin[1]_net_1 ), .Y(\n_din[5] ));
    crc16_2 UCRC3 (.crc3({\crc3[14] , \crc3[13] , \crc3[12] , 
        \crc3[11] , \crc3[10] , \crc3[9] , \crc3[8] , \crc3[7] , 
        \crc3[6] , \crc3[5] , \crc3[4] , \crc3[3] , \crc3[2] , 
        \crc3[1] , \crc3[0] }), .bits_0(\bits[3]_net_1 ), .crc_en(
        crc_en_net_1), .sdclk_n_1(sdclk_n_1), .crc_clr_i(crc_clr_i));
    CFG4 #( .INIT(16'h80BF) )  \n_bits_15_i_m4[3]  (.A(\crc3[10] ), .B(
        \i[2]_net_1 ), .C(\i[0]_net_1 ), .D(
        \n_bits_15_i_m4_1[3]_net_1 ), .Y(N_3791));
    CFG3 #( .INIT(8'hFE) )  data_bus_busy_RNO_0 (.A(\state[5]_net_1 ), 
        .B(\state[1]_net_1 ), .C(\state[0]_net_1 ), .Y(N_383_i));
    CFG2 #( .INIT(4'h4) )  \n_din[11]  (.A(\state[0]_net_1 ), .B(
        \odin[7]_net_1 ), .Y(\n_din[11]_net_1 ));
    CFG3 #( .INIT(8'h8D) )  n_wen7_RNISL0R (.A(\state[2]_net_1 ), .B(
        n_wen7_net_1), .C(N_386_i), .Y(un1_n_data_bus_busy8_2_i));
    CFG3 #( .INIT(8'h12) )  \n_blkn[0]  (.A(\blkn[0]_net_1 ), .B(
        \state[0]_net_1 ), .C(un1_n_blkn_0_sqmuxa_net_1), .Y(
        \n_blkn[0]_net_1 ));
    CFG3 #( .INIT(8'h12) )  \blkn_RNO[2]  (.A(\blkn[2]_net_1 ), .B(
        \state[0]_net_1 ), .C(CO1), .Y(N_3770_i));
    CFG4 #( .INIT(16'hCECC) )  \state_ns_0[1]  (.A(\state[3]_net_1 ), 
        .B(\state_ns_0_0[1]_net_1 ), .C(N_702), .D(n_dq8), .Y(
        \state_ns[1] ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_10_0_0_wmux[3]  (.A(
        \i[0]_net_1 ), .B(\i[3]_net_1 ), .C(\crc3[13] ), .D(\crc3[12] )
        , .FCI(VCC_net_1), .S(), .Y(\n_bits_10_0_0_y0[3] ), .FCO(
        \n_bits_10_0_0_co0[3] ));
    ARI1 #( .INIT(20'h0F588) )  \bits_ldmx_4_1_0_wmux_0[0]  (.A(
        \bits_ldmx_4_1_0_y0[0] ), .B(\bits_en[0]_net_1 ), .C(
        \bits_ldmx_2[0]_net_1 ), .D(N_3934_i), .FCI(
        \bits_ldmx_4_1_0_co0[0] ), .S(), .Y(
        \bits_ldmx_4_1_0_wmux_0_Y[0] ), .FCO());
    CFG4 #( .INIT(16'h1BB0) )  \n_i_0_iv_0[4]  (.A(n_i_sn_N_7_mux), .B(
        \n_i_0_iv_0_1[4]_net_1 ), .C(\i[4]_net_1 ), .D(un48_n_i_c4), 
        .Y(\n_i_0_iv_0[4]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \state_ns_0_a2_0[5]  (.A(N_137), .B(
        \state[5]_net_1 ), .C(un1_i_4lt4), .D(
        \state_ns_0_a2_0_1_1_a2_1[5]_net_1 ), .Y(N_729));
    CFG4 #( .INIT(16'hEA40) )  \i_lm_0[7]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(un1_state_21_i), .C(
        \i[7]_net_1 ), .D(\i_s[7] ), .Y(\i_lm[7] ));
    CFG3 #( .INIT(8'h84) )  \n_i_iv_0_a2_s[0]  (.A(\i[0]_net_1 ), .B(
        \state[4]_net_1 ), .C(status_0), .Y(n_i_iv_0_a2_out));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[6]  (.A(\state[0]_net_1 ), .B(
        \odin[2]_net_1 ), .Y(N_70_i));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    SLE \state[2]  (.D(N_687_i), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[2]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \n_dq_0[2]  (.A(\data0[2]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\n_dq_0[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[21]  (.A(\state[0]_net_1 ), .B(
        \odin[17]_net_1 ), .Y(\n_din[21] ));
    SLE \bits[3]  (.D(\bits_ldmx[3]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_data_out_en_3_sqmuxa_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\bits[3]_net_1 ));
    CFG4 #( .INIT(16'hFEF0) )  un1_state_21_0_0_1 (.A(\dq[2]_net_1 ), 
        .B(\dq[3]_net_1 ), .C(\state[4]_net_1 ), .D(\state[1]_net_1 ), 
        .Y(un1_state_21_0_0_1_net_1));
    CFG4 #( .INIT(16'hECA0) )  \state_ns_0_0[1]  (.A(sd_write_start), 
        .B(\state[1]_net_1 ), .C(\state[0]_net_1 ), .D(N_700), .Y(
        \state_ns_0_0[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_s[9]  (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[8]_net_1 ), .S(\i_s[9]_net_1 ), .Y(), .FCO());
    SLE is_last_data_inst_1 (.D(n_is_last_data_iv_i), .CLK(sdclk_n_1), 
        .EN(N_384_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(is_last_data));
    CFG3 #( .INIT(8'h80) )  n_is_last_data_iv_0_a3 (.A(n_dq8), .B(
        \state[3]_net_1 ), .C(N_702_i), .Y(N_3819));
    SLE \state[1]  (.D(\state_ns[1] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[8]  (.A(din[4]), .B(
        \odin[4]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(\n_AX[8] )
        );
    SLE \AX[1]  (.D(N_3768_i), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[1]));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    SLE \i[5]  (.D(\i_lm[5] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    CFG4 #( .INIT(16'h1011) )  n_data_out_2_sqmuxa_2_RNIPS4B1 (.A(
        \state[1]_net_1 ), .B(\state[2]_net_1 ), .C(N_702_i), .D(
        n_data_out_2_sqmuxa_2_net_1), .Y(un1_state_9_i));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[30]  (.A(din[26]), .B(
        \odin[26]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[30] ));
    CFG4 #( .INIT(16'h8000) )  n_is_last_data6 (.A(\i[0]_net_1 ), .B(
        \i[2]_net_1 ), .C(n_is_last_data6_4_net_1), .D(
        n_is_last_data6_3_0_net_1), .Y(n_is_last_data6_net_1));
    CFG4 #( .INIT(16'hEA40) )  \i_lm_0[9]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(un1_state_21_i), .C(
        \i[9]_net_1 ), .D(\i_s[9]_net_1 ), .Y(\i_lm[9] ));
    SLE \i[8]  (.D(\i_lm[8] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    SLE \data0[0]  (.D(sd_data_in[0]), .CLK(sdclk_n_i), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\data0[0]_net_1 ));
    SLE \AX[16]  (.D(\n_AX[16] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[16]));
    SLE \AX[5]  (.D(\n_AX[5] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[5]));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_13_i_m3_0_0_wmux_0[3]  (.A(
        \n_bits_13_i_m3_0_0_y0[3] ), .B(\i[0]_net_1 ), .C(\crc3[6] ), 
        .D(\crc3[2] ), .FCI(\n_bits_13_i_m3_0_0_co0[3] ), .S(), .Y(
        N_3778), .FCO());
    CFG3 #( .INIT(8'hBA) )  \state_ns_i_0[6]  (.A(N_731), .B(
        \state[7]_net_1 ), .C(N_386_i), .Y(\state_ns_i_0[6]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[17]  (.A(\state[0]_net_1 ), .B(
        \odin[13]_net_1 ), .Y(\n_din[17] ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[13]  (.A(din[9]), .B(
        \odin[9]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[13] ));
    CFG4 #( .INIT(16'hF4E4) )  \n_i_0_iv_0[5]  (.A(n_i_sn_N_7_mux), .B(
        n_i_0_iv_0_a2_1_out), .C(\i[5]_net_1 ), .D(\state[4]_net_1 ), 
        .Y(\n_i_0_iv_0[5]_net_1 ));
    CFG3 #( .INIT(8'h53) )  \bits_ldmx_1[3]  (.A(N_818), .B(
        \bits[3]_net_1 ), .C(\bits_en[0]_net_1 ), .Y(
        \bits_ldmx_1[3]_net_1 ));
    CFG4 #( .INIT(16'hB888) )  \i_lm_0[5]  (.A(\i_s[5] ), .B(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .C(un1_state_21_i), .D(
        \n_i_0_iv_0[5]_net_1 ), .Y(\i_lm[5] ));
    CFG2 #( .INIT(4'h4) )  \odin_RNO[7]  (.A(\state[0]_net_1 ), .B(
        \odin[3]_net_1 ), .Y(N_68_i));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(\i_cry[5]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \un18_0_a2[2]  (.A(\state[7]_net_1 ), .B(
        \state[4]_net_1 ), .C(N_386_i), .Y(N_378));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_12_i_m2_0_0_wmux[1]  (.A(
        \i[3]_net_1 ), .B(\i[0]_net_1 ), .C(\crc1[9] ), .D(\crc1[1] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_12_i_m2_0_0_y0[1] ), .FCO(
        \n_bits_12_i_m2_0_0_co0[1] ));
    ARI1 #( .INIT(20'h4AA00) )  i_s_417 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(i_s_417_FCO));
    CFG2 #( .INIT(4'h4) )  \n_din[15]  (.A(\state[0]_net_1 ), .B(
        \odin[11]_net_1 ), .Y(\n_din[15]_net_1 ));
    CFG4 #( .INIT(16'h1101) )  \n_bits_16_i_0_RNIN5V01[0]  (.A(
        \n_bits_16_i_0[0]_net_1 ), .B(\n_bits_16_i_1[0]_net_1 ), .C(
        un1_i_4lt4), .D(N_3941), .Y(N_3934_i));
    CFG3 #( .INIT(8'h80) )  \un1_blkn_1.CO1  (.A(\blkn[0]_net_1 ), .B(
        un1_n_blkn_0_sqmuxa_net_1), .C(\blkn[1]_net_1 ), .Y(CO1));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[12]  (.A(din[8]), .B(
        \odin[8]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[12] ));
    CFG4 #( .INIT(16'hFFFE) )  \state_ns_0_o4[1]  (.A(\dq[3]_net_1 ), 
        .B(\dq[2]_net_1 ), .C(\dq[1]_net_1 ), .D(\dq[0]_net_1 ), .Y(
        N_700));
    CFG2 #( .INIT(4'h7) )  \state_ns_0_o4_1[3]  (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .Y(\state_ns_0_o4_1[3]_net_1 ));
    SLE \AX[26]  (.D(\n_AX[26] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[26]));
    CFG3 #( .INIT(8'h8E) )  \n_dq8_1.CO2  (.A(CO2_1), .B(
        total_blocks[2]), .C(\blkn[2]_net_1 ), .Y(CO2));
    CFG4 #( .INIT(16'h7222) )  \i_lm_0[0]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(\i[0]_net_1 ), .C(
        un1_state_21_i), .D(\i_lm_0_1_0[0]_net_1 ), .Y(\i_lm[0] ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[10]  (.A(din[6]), .B(
        \odin[6]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[10] ));
    CFG2 #( .INIT(4'h1) )  \i_RNI53PC[8]  (.A(\i[8]_net_1 ), .B(
        \i[9]_net_1 ), .Y(N_137));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_10_i_m2_0_0_wmux_0[1]  (.A(
        \n_bits_10_i_m2_0_0_y0[1] ), .B(\i[3]_net_1 ), .C(\crc1[5] ), 
        .D(\crc1[4] ), .FCI(\n_bits_10_i_m2_0_0_co0[1] ), .S(), .Y(
        N_3947), .FCO());
    SLE \i[3]  (.D(\i_lm[3] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    CFG2 #( .INIT(4'hE) )  data_bus_busy_RNO (.A(\state[1]_net_1 ), .B(
        \state[5]_net_1 ), .Y(N_387_i));
    CFG4 #( .INIT(16'hD888) )  \i_lm_0[4]  (.A(
        \state_ns_0_a2_0_RNI7N2R[5]_net_1 ), .B(\i_s[4] ), .C(
        un1_state_21_i), .D(\n_i_0_iv_0[4]_net_1 ), .Y(\i_lm[4] ));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[4]  (.A(\state[0]_net_1 ), .B(
        \odin[0]_net_1 ), .Y(\n_din[4] ));
    CFG2 #( .INIT(4'h4) )  \n_din[20]  (.A(\state[0]_net_1 ), .B(
        \odin[16]_net_1 ), .Y(\n_din[20]_net_1 ));
    SLE \odin[4]  (.D(\n_din[4] ), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[4]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[29]  (.A(din[25]), .B(
        \odin[25]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[29] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[8]  (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[7]_net_1 ), .S(\i_s[8] ), .Y(), .FCO(\i_cry[8]_net_1 ));
    CFG2 #( .INIT(4'h4) )  crc_clr_RNO_1 (.A(N_135), .B(
        \state[7]_net_1 ), .Y(N_76_i));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[31]  (.A(din[27]), .B(
        \odin[27]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[31] ));
    SLE \AX[8]  (.D(\n_AX[8] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[8]));
    CFG3 #( .INIT(8'h01) )  un1_state_18_1 (.A(\state[4]_net_1 ), .B(
        \state[0]_net_1 ), .C(\state[1]_net_1 ), .Y(
        un1_state_18_1_net_1));
    CFG3 #( .INIT(8'h53) )  \bits_ldmx_1[1]  (.A(N_816), .B(
        \bits[1]_net_1 ), .C(\bits_en[0]_net_1 ), .Y(
        \bits_ldmx_1[1]_net_1 ));
    SLE \i[1]  (.D(\i_lm[1] ), .CLK(sdclk_n_1), .EN(N_3446_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_din_0_a2[16]  (.A(\state[0]_net_1 ), .B(
        \odin[12]_net_1 ), .Y(\n_din[16] ));
    CFG4 #( .INIT(16'h0051) )  \state_ns_0_a2_RNITNV31[4]  (.A(
        \state[2]_net_1 ), .B(\state[3]_net_1 ), .C(n_data_out6_net_1), 
        .D(N_726), .Y(un1_state_6_i));
    CFG4 #( .INIT(16'hA808) )  n_data_out_1_sqmuxa_1 (.A(
        \state[3]_net_1 ), .B(\i[1]_net_1 ), .C(\i[2]_net_1 ), .D(
        \i[0]_net_1 ), .Y(n_data_out_1_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'h6A00) )  \n_i_0_iv_0_a2_1_s[5]  (.A(\i[5]_net_1 )
        , .B(\i[4]_net_1 ), .C(un48_n_i_c4), .D(
        \n_i_iv_0_a2_2_0[0]_net_1 ), .Y(n_i_0_iv_0_a2_1_out));
    SLE \data0[2]  (.D(sd_data_in[2]), .CLK(sdclk_n_i), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\data0[2]_net_1 ));
    SLE \AX[2]  (.D(\n_AX[2] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[2]));
    CFG3 #( .INIT(8'hB8) )  \n_bits_9[1]  (.A(din[29]), .B(
        \state[6]_net_1 ), .C(n_bits_17_sqmuxa), .Y(N_787));
    CFG3 #( .INIT(8'hE4) )  \n_bits_16_bm[1]  (.A(\i[2]_net_1 ), .B(
        N_3947), .C(N_3945), .Y(\n_bits_16_bm[1]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_10_i_m2_0_0_wmux[1]  (.A(
        \i[0]_net_1 ), .B(\i[3]_net_1 ), .C(\crc1[13] ), .D(\crc1[12] )
        , .FCI(VCC_net_1), .S(), .Y(\n_bits_10_i_m2_0_0_y0[1] ), .FCO(
        \n_bits_10_i_m2_0_0_co0[1] ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[24]  (.A(din[20]), .B(
        \odin[20]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[24] ));
    CFG4 #( .INIT(16'h33BA) )  \i_lm_0_1_0[0]  (.A(n_i_iv_0_a2_out), 
        .B(\i[0]_net_1 ), .C(\n_i_iv_0_a2_2_0[0]_net_1 ), .D(
        n_i_sn_N_7_mux), .Y(\i_lm_0_1_0[0]_net_1 ));
    SLE \odin[22]  (.D(N_64_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[22]_net_1 ));
    SLE \odin[12]  (.D(\n_din[12] ), .CLK(sdclk_n_1), .EN(N_388_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\odin[12]_net_1 ));
    CFG4 #( .INIT(16'h80BF) )  \n_bits_16_i_m2_1[0]  (.A(\crc0[12] ), 
        .B(\i[1]_net_1 ), .C(\i[0]_net_1 ), .D(
        \n_bits_16_i_m2_1_1[0]_net_1 ), .Y(N_3941));
    SLE \data_out[0]  (.D(\n_data_out_iv_i_0[0]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_9_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sd_data_out[0]));
    SLE \blkn[1]  (.D(\n_blkn[1]_net_1 ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \blkn[1]_net_1 ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv_0[21]  (.A(din[17]), .B(
        \odin[17]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[21] ));
    SLE \odin[6]  (.D(N_70_i), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[6]_net_1 ));
    ARI1 #( .INIT(20'h0FA44) )  \n_bits_12_0_0_wmux[2]  (.A(
        \i[3]_net_1 ), .B(\i[0]_net_1 ), .C(\crc2[9] ), .D(\crc2[1] ), 
        .FCI(VCC_net_1), .S(), .Y(\n_bits_12_0_0_y0[2] ), .FCO(
        \n_bits_12_0_0_co0[2] ));
    CFG4 #( .INIT(16'hCE0A) )  \n_AX_iv[20]  (.A(din[16]), .B(
        \odin[16]_net_1 ), .C(N_78), .D(\state[2]_net_1 ), .Y(
        \n_AX[20] ));
    CFG4 #( .INIT(16'h0031) )  is_last_data_RNO (.A(\state[2]_net_1 ), 
        .B(\state[0]_net_1 ), .C(n_is_last_data6_net_1), .D(N_3819), 
        .Y(n_is_last_data_iv_i));
    CFG3 #( .INIT(8'h80) )  n_wen7 (.A(\i[2]_net_1 ), .B(\i[0]_net_1 ), 
        .C(\i[1]_net_1 ), .Y(n_wen7_net_1));
    ARI1 #( .INIT(20'h0F588) )  \n_bits_13_i_m3_0_0_wmux_0[1]  (.A(
        \n_bits_13_i_m3_0_0_y0[1] ), .B(\i[0]_net_1 ), .C(\crc1[6] ), 
        .D(\crc1[2] ), .FCI(\n_bits_13_i_m3_0_0_co0[1] ), .S(), .Y(
        N_3780), .FCO());
    ARI1 #( .INIT(20'h0F588) )  \n_bits_13_i_m2_0_0_wmux_0[0]  (.A(
        \n_bits_13_i_m2_0_0_y0[0] ), .B(\i[0]_net_1 ), .C(\crc0[6] ), 
        .D(\crc0[2] ), .FCI(\n_bits_13_i_m2_0_0_co0[0] ), .S(), .Y(
        N_3944), .FCO());
    SLE \AX[7]  (.D(\n_AX[7] ), .CLK(sdclk_n_1), .EN(
        un1_n_data_bus_busy8_2_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(din[7]));
    CFG2 #( .INIT(4'h4) )  \n_din[19]  (.A(\state[0]_net_1 ), .B(
        \odin[15]_net_1 ), .Y(\n_din[19]_net_1 ));
    SLE \odin[5]  (.D(\n_din[5] ), .CLK(sdclk_n_1), .EN(N_388_i), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\odin[5]_net_1 ));
    
endmodule


module sdtop(
       test_0_HADDR,
       test_0_HWDATA,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0,
       sd_data_in,
       sd_data_out,
       test_0_HTRANS_0,
       test_0_HADDR_i_0,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       test_0_HWRITE,
       spdif_tx_c,
       olrck_o,
       reset_n_i_2,
       reset_n_i_i_2,
       reset_n_i_3,
       reset_n_i_i_1,
       reset_n_i_1,
       reset_n_i_i_0,
       reset_n_i_0,
       mclk_1,
       reset_n_i_i,
       sd_data_out_en_i_i,
       data_out_en_ret_fast_i,
       odata_o,
       obck_o,
       cmd_in,
       sdclk_n_i,
       cmd_out,
       spdif_en_c,
       en49_c,
       en45_c,
       sdclk_n_1,
       u8_sb_0_HPMS_READY,
       cmd_out_en_i_i
    );
output [16:2] test_0_HADDR;
output [31:0] test_0_HWDATA;
input  [31:0] u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0;
input  [3:0] sd_data_in;
output [3:0] sd_data_out;
output test_0_HTRANS_0;
output test_0_HADDR_i_0;
input  u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
output test_0_HWRITE;
output spdif_tx_c;
output olrck_o;
output reset_n_i_2;
input  reset_n_i_i_2;
output reset_n_i_3;
input  reset_n_i_i_1;
output reset_n_i_1;
input  reset_n_i_i_0;
output reset_n_i_0;
input  mclk_1;
input  reset_n_i_i;
output sd_data_out_en_i_i;
output data_out_en_ret_fast_i;
output odata_o;
output obck_o;
input  cmd_in;
input  sdclk_n_i;
output cmd_out;
output spdif_en_c;
output en49_c;
output en45_c;
input  sdclk_n_1;
input  u8_sb_0_HPMS_READY;
output cmd_out_en_i_i;

    wire reset_n_i_0_RNIOUJE_net_1, reset_n_i_0_0, cmd_out_en_i, N_845, 
        N_845_i, dsd_clkr_i_i, N_4047_i, crc_clr_net_1, crc_clr_i, 
        \total_blocks[3]_net_1 , VCC_net_1, \n_total_blocks[3]_net_1 , 
        N_152_i, GND_net_1, \cccr_func_sel[0]_net_1 , N_77_i, un87_i, 
        \cccr_func_sel[1]_net_1 , N_3651_i, \cccr_func_sel[2]_net_1 , 
        N_3650_i, \cccr_func_sel[3]_net_1 , N_3649_i, \ind[0]_net_1 , 
        ind_389_net_1, \ind[1]_net_1 , ind_390_net_1, \ind[2]_net_1 , 
        ind_391_net_1, \ind[3]_net_1 , ind_392_net_1, \ind[4]_net_1 , 
        ind_393_net_1, \ind[5]_net_1 , ind_394_net_1, 
        \total_blocks[0]_net_1 , \n_total_blocks[0]_net_1 , 
        \total_blocks[1]_net_1 , \n_total_blocks[1]_net_1 , 
        \total_blocks[2]_net_1 , \n_total_blocks[2]_net_1 , 
        \sound_card_ctrl[5]_net_1 , N_3648_i, un105_i_0_net_1, 
        \sound_card_ctrl[6]_net_1 , N_3647_i, 
        \sound_card_ctrl[7]_net_1 , N_3646_i, 
        \sound_card_ctrl[0]_net_1 , un102_i_0_net_1, 
        \sound_card_ctrl[1]_net_1 , \sound_card_ctrl[2]_net_1 , 
        \arg[0]_net_1 , n_sound_card_ctrl_1_sqmuxa_1, \arg[1]_net_1 , 
        \response[25]_net_1 , \n_response_1[25] , un1_state_11_i, 
        \response[26]_net_1 , \n_response_1[26] , \response[27]_net_1 , 
        \n_response_1[27] , \response[28]_net_1 , \n_response_1[28] , 
        \response[29]_net_1 , \n_response_1[29] , \response[30]_net_1 , 
        \n_response_1[30] , \response[31]_net_1 , \n_response_1[31] , 
        \response[32]_net_1 , \n_response_1[32] , \response[33]_net_1 , 
        \n_response_1[33] , \response[34]_net_1 , 
        \n_response_1_1_iv_i[34] , \response[35]_net_1 , 
        \n_response_1[35] , \response[36]_net_1 , 
        \n_response_1_1_iv_i[36] , \response[37]_net_1 , 
        \n_response_1_1_iv_i[37] , \response[38]_net_1 , 
        \n_response_1[38] , \response[39]_net_1 , \n_response_1[39] , 
        \response[12]_net_1 , \n_response_1_0_iv_i[12] , 
        \response[13]_net_1 , \n_response_1[13] , \response[14]_net_1 , 
        \n_response_1[14] , \response[15]_net_1 , \n_response_1[15] , 
        \response[16]_net_1 , \n_response_1[16] , \response[17]_net_1 , 
        \n_response_1[17] , \response[18]_net_1 , \n_response_1[18] , 
        \response[19]_net_1 , \n_response_1[19] , \response[20]_net_1 , 
        \n_response_1[20] , \response[21]_net_1 , \n_response_1[21] , 
        \response[22]_net_1 , \n_response_1[22] , \response[23]_net_1 , 
        \n_response_1[23] , \response[24]_net_1 , \n_response_1[24] , 
        \arg[27]_net_1 , arg_372_net_1, \arg[28]_net_1 , arg_373_net_1, 
        \arg[29]_net_1 , arg_374_net_1, \arg[30]_net_1 , arg_375_net_1, 
        \arg[31]_net_1 , arg_376_net_1, \response[0]_net_1 , 
        \n_response_1[0] , \response[2]_net_1 , \n_response_1[2] , 
        \response[3]_net_1 , \n_response_1[3] , \response[4]_net_1 , 
        \n_response_1[4] , \response[5]_net_1 , \n_response_1[5] , 
        \response[6]_net_1 , \n_response_1[6] , \response[7]_net_1 , 
        \n_response_1[7] , \response[8]_net_1 , \n_response_1[8] , 
        \arg[12]_net_1 , arg_357_net_1, \arg[13]_net_1 , arg_358_net_1, 
        \arg[14]_net_1 , arg_359_net_1, \arg[15]_net_1 , arg_360_net_1, 
        \arg[16]_net_1 , arg_361_net_1, \arg[17]_net_1 , arg_362_net_1, 
        \arg[18]_net_1 , arg_363_net_1, \arg[19]_net_1 , arg_364_net_1, 
        \arg[20]_net_1 , arg_365_net_1, \arg[21]_net_1 , arg_366_net_1, 
        \arg[22]_net_1 , arg_367_net_1, \arg[23]_net_1 , arg_368_net_1, 
        \arg[24]_net_1 , arg_369_net_1, \arg[25]_net_1 , arg_370_net_1, 
        \arg[26]_net_1 , arg_371_net_1, N_342, un77, \n_arg[1]_net_1 , 
        \arg[2]_net_1 , \n_arg[2]_net_1 , \arg[3]_net_1 , 
        \n_arg[3]_net_1 , \arg[4]_net_1 , \n_arg[4]_net_1 , 
        \arg[5]_net_1 , \n_arg[5]_net_1 , \arg[6]_net_1 , 
        \n_arg[6]_net_1 , \arg[7]_net_1 , \n_arg[7]_net_1 , 
        \arg[8]_net_1 , \n_arg[8] , \arg[9]_net_1 , arg_354_net_1, 
        \arg[10]_net_1 , arg_355_net_1, \arg[11]_net_1 , arg_356_net_1, 
        sd_read_start_net_1, \state[10]_net_1 , un107_i, 
        \state[2]_net_1 , N_144, in_cmd_net_1, \state[1]_net_1 , 
        un97_i_a6_net_1, n_spdif_en_1_sqmuxa, cmd_q2_net_1, N_341_i, 
        un103_i_a6_net_1, n_cmd_out_iv_i, un95_i_0_net_1, no_crc_net_1, 
        no_crc_397_net_1, crc_en_net_1, N_3522_i, N_1699, 
        sd_write_start_net_1, N_2938_i, un101_i, cccr_reset_net_1, 
        cccr_reset_388_net_1, cmd_q_net_1, n_cmd_q_net_1, 
        cccr_cd_disable_net_1, n_cccr_cd_disable_1_sqmuxa_net_1, 
        bit_net_1, \state[3]_net_1 , \state_ns[3] , \state[4]_net_1 , 
        N_2223_i, \state[5]_net_1 , N_4042_i, \state[6]_net_1 , 
        \state_ns[6] , \state[7]_net_1 , \state_ns[7] , 
        \state[8]_net_1 , \state_ns[8] , \state[9]_net_1 , N_2163_i, 
        \state_ns[10] , \state[11]_net_1 , N_2166_i, \state[12]_net_1 , 
        N_2168_i, \state[0]_net_1 , N_154_i, N_2153_i, \state_ns[2] , 
        \bus_state[0]_net_1 , \bus_state_ns[0] , \bus_state[1]_net_1 , 
        \bus_state_ns[1] , \bus_state[2]_net_1 , \bus_state_ns[2] , 
        \bus_state[3]_net_1 , \bus_state_ns[3] , \bus_state[4]_net_1 , 
        N_2263_i, cmd0_net_1, in_bck_1, start_dsd_tx_net_1, dsd_clk_1, 
        dop_start, start_pcm_tx_net_1, start_pcm_tx_2, \i[6]_net_1 , 
        \i_lm[6] , \i[7]_net_1 , \i_lm[7] , 
        \buffer_under_run[0]_net_1 , \buffer_under_run_s[0] , 
        buffer_under_rune, \buffer_under_run[1]_net_1 , 
        \buffer_under_run_s[1] , \buffer_under_run[2]_net_1 , 
        \buffer_under_run_s[2] , \buffer_under_run[3]_net_1 , 
        \buffer_under_run_s[3] , \buffer_under_run[4]_net_1 , 
        \buffer_under_run_s[4] , \buffer_under_run[5]_net_1 , 
        \buffer_under_run_s[5] , \buffer_under_run[6]_net_1 , 
        \buffer_under_run_s[6] , \buffer_under_run[7]_net_1 , 
        \buffer_under_run_s[7] , cmd_out_en_i_reti, un96_i_0_net_1, 
        N_2431_reto, N_2431, N_3732_reto, N_3732, \i_reto[0] , \i[0] , 
        \i_s_reto[0] , \i_s[0] , \n_response_1_0_iv_2_reto[1] , 
        \n_response_1_0_iv_2[1]_net_1 , \n_response_123_m_reto[1] , 
        \n_response_123_m[1]_net_1 , \n_response_360_reto[1] , 
        \n_response_360[1] , \state_reto[9] , 
        \n_response_1_0_iv_0_reto[11] , 
        \n_response_1_0_iv_0[11]_net_1 , \n_response_406_m_reto[11] , 
        \n_response_406_m[11] , \n_response_cnst_1_m_reto[9] , 
        \n_response_cnst_1_m[9] , N_3595_reto, N_3595, 
        \n_response_cnst_1_m_reto_0[9] , \response_reto[10] , 
        \response[10] , \response_m_0_reto[9] , \response_m_0[9] , 
        N_845_reto, \n_response_1_0_iv_0_reto[9] , 
        \n_response_1_0_iv_0[9]_net_1 , 
        \n_response_cnst_1_m_reto_1[9] , \response_reto[8] , 
        N_3732_reto_0, N_3737_reto, N_3737, N_3738_reto, N_3738, 
        \i_s_reto[3] , \i_s[3] , N_73_reto, N_73, N_74_reto, N_74, 
        N_3732_reto_1, \i_s_reto[2] , \i_s[2] , N_3732_reto_2, 
        \i_s_reto[1] , \i_s[1] , \n_i_reto[1] , \n_i[1] , \i[5]_net_1 , 
        \i_lm[5] , \i[4]_net_1 , \i_lm[4] , i_cry_cy, N_1407_i, N_3762, 
        n_state_3_sqmuxa_0_a4_i_1_0, \i_cry[0]_net_1 , \i_0[0] , 
        \i_qxu[0]_net_1 , \i_cry[1]_net_1 , \i_cry[2]_net_1 , \i_0[2] , 
        \i_qxu[2]_net_1 , \i_cry[3]_net_1 , \i_0[3] , \i_qxu[3]_net_1 , 
        \i_cry[4]_net_1 , \i_s[4] , 
        n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1, un1_i_3, 
        \i_cry[5]_net_1 , \i_s[5] , \i_s[7]_net_1 , \i_cry[6]_net_1 , 
        \i_s[6] , buffer_under_run_cry_cy, \buffer_under_run_cry[0] , 
        \buffer_under_run_cry[1] , \buffer_under_run_cry[2] , 
        \buffer_under_run_cry[3] , \buffer_under_run_cry[4] , 
        \buffer_under_run_cry[5] , \buffer_under_run_cry[6] , N_702, 
        \n_response_49_4_1[7] , n_state_0_sqmuxa_0_a6_0_a3_1_net_1, 
        n_state_0_sqmuxa, un1_arg_13_i_i_a2_0_13_2, 
        un1_arg_13_i_i_a2_0_13_4, N_1697, \n_response_360_1[0]_net_1 , 
        N_709, \n_response_360_m[0] , N_213_i, N_3724, N_1696_i, 
        N_979_1, N_1684, un101_2_net_1, 
        \n_response_1_0_iv_0_m2_6_1_1[5] , 
        \n_response_1_0_iv_0_m2_6_1[5] , N_12, N_55, N_66_mux, N_3572, 
        \n_response_360_4_1_1[1] , \response[1] , m31_s, 
        \n_response_360_4_1[1] , N_4044_i, N_4043_i, \n_i[4] , N_69, 
        N_3534, \i[1] , \i[2] , \i[3] , \n_response_360_1_0[3]_net_1 , 
        n_response_360_0_net_1, \n_response_360[3]_net_1 , N_334, 
        m42_0_2, \n_response_360_1_0[7]_net_1 , 
        \n_response_360[7]_net_1 , N_60, \n_response_360_1_0[2]_net_1 , 
        \n_response_360[2]_net_1 , i4_mux_1, N_2221, 
        \state_ns_0_4[3]_net_1 , \state_ns_0_1_0[3]_net_1 , N_2218, 
        \state_ns_0_a3_4_1[3]_net_1 , N_2222_1_0, N_970, 
        n_cmd_out_iv_0_a2_1_2, N_147, n_cmd_out_iv_0_a2_7_1_0_net_1, 
        \bus_state_ns_0_1[3]_net_1 , \bus_state_ns_0_0[3]_net_1 , 
        N_1686_i, N_2266, N_4043_i_1, N_243, N_634_1, m59_1_1, N_1163, 
        N_11, N_2263_i_1, N_3666, N_1386_i, n_state42, N_4044_i_1, 
        \n_response_49_1_1[6]_net_1 , \n_response_36[6]_net_1 , 
        \n_response_49[6]_net_1 , n_response_49_4_net_1, N_2537, 
        \n_response_49_1[2]_net_1 , \n_response_49[2]_net_1 , N_1166, 
        N_706, n_response_49_8_net_1, N_2538, 
        \n_response_49_1[3]_net_1 , \n_response_49[3]_net_1 , 
        n_response_6_sqmuxa_1_net_1, N_4040, n_response_6_sqmuxa_net_1, 
        \n_response_36_1_1[6]_net_1 , \status[6] , N_1164, N_49, 
        m50_1_0, \n_response_cnst_4[4] , m48_1_1, 
        n_response_4_sqmuxa_i_1, N_4, m54_0_1, m54_0, 
        \n_response_49_0[7]_net_1 , \n_response_49[7] , 
        \n_response_49_4_1_0[1] , \n_response_36[1]_net_1 , 
        \n_response_49_4_1_1[1] , \n_response_49[1] , 
        \n_response_360_0[0]_net_1 , m17_s, m17_d_s, m17_d_d, i4_mux_0, 
        \status[7] , N_2541, N_4038_i, N_702_1, N_3634_2, N_3634, 
        un107_0_0_net_1, N_3528, N_244, un103_i_a6_0_net_1, 
        n_response_4_sqmuxa_0_a3_0_net_1, m16_1, N_181, 
        \n_response_159_m_xx_0[0]_net_1 , un1_arg_0_1_0_0, N_3641, 
        m42_0_a3_0, \state_ns_0_a2_0_a2_i_o3_0[3]_net_1 , 
        n_state_3_sqmuxa_0_a4_i_c, N_401, N_180, N_1166_i_2, 
        \response[9] , N_357_i, \response_i_m[1] , N_3736_1, N_3694, 
        N_3713, N_174, un1_arg_12_7, N_3589_i, N_2175_i_1, N_612, 
        n_response_3_sqmuxa_1, N_372, N_685_3, N_4039, N_4053, N_4054, 
        N_408, N_96_i, un72, un1_arg_12_12_net_1, N_355, N_276, 
        N_1387_i, N_374, n_state13_net_1, N_204, N_3592, use_dsd, 
        odata2, odata1, N_1165, N_4049, n_response_0_sqmuxa_1_net_1, 
        \n_response_1_0_iv_0[3]_net_1 , n_state_3_sqmuxa_0_a4_i_0_1, 
        \n_response_1_0_iv_0[1]_net_1 , \n_response_1_0_iv_0[7]_net_1 , 
        \n_response_1_0_iv_0[2]_net_1 , \n_response_1_0_iv_0[6]_net_1 , 
        un1_state_11_2_net_1, data_bus_busy, 
        \bus_state_ns_0_a4_1_1[3]_net_1 , 
        \n_response_1_0_iv_0_a3_5_1[4]_net_1 , un1_arg_15_1_net_1, 
        un1_arg_15_0_net_1, n_response_1_sqmuxa_6_1, 
        un1_arg_12_5_net_1, un1_arg_12_4_net_1, un1_arg_12_3_0, 
        \state_ns_0_a3_0_a2_i_1[5]_net_1 , 
        buffer_under_runlde_0_a6_0_1, un1_arg_13_i_i_a2_0_12_4, 
        un1_arg_13_i_i_a2_0_12_3, un1_arg_13_i_i_a2_0_13_1, 
        \state_ns_0_a3_0_a2_4_a3_1[10]_net_1 , 
        \state_ns_0_a3_0_a2_0_a3_1[6]_net_1 , 
        \state_ns_0_a3_3_0_a3_1[3]_net_1 , \state_ns_0_i_a2_0_0[0] , 
        n_state_2_sqmuxa_0_a6_a0_0, \state_ns_0_a3_2_0_0[3] , 
        n_state42_0_a2_0_a3_0_net_1, \state_ns_0_a3_0_0[7]_net_1 , 
        n_cmd_out_iv_0_a2_1_1_net_1, 
        n_cmd_out_en_1_sqmuxa_0_0_a3_0_2_1, N_678, cccr_cd_disable_m, 
        un1_arg_12_21_net_1, N_1016_3, N_3538, n_response_1_sqmuxa_2, 
        N_1061_1_0, N_221, N_318_4, N_290, N_795, N_289, 
        un1_buffer_under_runlt5, N_3579, \n_response_159_m[3]_net_1 , 
        \n_response_123_m[6]_net_1 , N_2222_10, N_967, N_1060, N_3747, 
        N_1013_3, N_1014_3, N_3692, N_1062_1_0, 
        \n_response_159_m_xx[1]_net_1 , un1_arg_12_22_0_net_1, 
        N_3736_4, un12_n_i_c3, \cccr_func_sel_m[3] , 
        \cccr_func_sel_m[2] , N_2265, N_2186, N_3696, N_3658, N_3630, 
        n_response_1_sqmuxa_net_1, N_300, \n_response_cnst_2[6] , 
        N_413, N_393, N_10, N_2721, N_229, N_3, N_659, \crc[1] , 
        \crc[0] , n_cmd_out_iv_0_a2_1_0_net_1, 
        \n_response_36[4]_net_1 , N_3574, N_3573, 
        n_state_3_sqmuxa_0_a4_i_0_2, \n_response_123_iv_0[0]_net_1 , 
        buffer_under_runlde_0_a6_5, \state_ns_0_i_o2_1[0]_net_1 , 
        \state_ns_0_i_o2_0[0]_net_1 , un1_n_response_3_sqmuxa_i_0, 
        un104_i_a6_1_net_1, n_response_5_sqmuxa_1_1_net_1, 
        \state_ns_0_a3_0_a2_i_2[5]_net_1 , un1_arg_1_1, un1_arg_0_0, 
        \state_ns_0_a3_0_0_a6_2[8]_net_1 , un95_i_a6_0_1_0_0_net_1, 
        n_cccr_reset_0_sqmuxa_1_0_net_1, 
        n_response_14_sqmuxa_1_tz_1_net_1, 
        n_cmd_out4_0_a2_0_a3_1_net_1, n_state_2_sqmuxa_0_a6_a0_net_1, 
        \state_ns_0_a2_3_1_a6_0_a2_3[0]_net_1 , \crc[6] , N_164, 
        N_2220, un1_buffer_under_runlt7, N_333, N_314, N_336, N_335, 
        N_313, \crc[4] , N_160, \crc[3] , N_163, N_318, N_3745, 
        n_state_1_sqmuxa, N_361, N_231, \n_response_159_m_xx[0]_net_1 , 
        un1_arg_12_22_net_1, \state_ns_0_i_o2_0_1[0]_net_1 , 
        n_response_16_sqmuxa_i_0_0_net_1, un12_n_i_c4, N_3654, 
        N_1061_2_0, N_2181, N_3524, \n_response_159_m[1] , 
        \n_response_159_m[2]_net_1 , \n_response_159[6]_net_1 , 
        n_sound_card_ctrl_2_sqmuxa, \response[11] , 
        \n_response_1_1_iv_0_0[37]_net_1 , 
        \n_response_1_0_iv_0_0[32]_net_1 , 
        \n_response_1_1_iv_0_0[36]_net_1 , 
        \n_response_1_1_iv_0_0[20]_net_1 , 
        \n_response_1_1_iv_0_0[31]_net_1 , 
        \n_response_1_1_iv_0_0[35]_net_1 , 
        \n_response_1_1_iv_0_0[17]_net_1 , 
        \n_response_1_1_iv_0_0[23]_net_1 , 
        \n_response_1_1_iv_0_0[28]_net_1 , 
        \n_response_1_1_iv_0_0[15]_net_1 , 
        \n_response_1_1_iv_0_0[18]_net_1 , 
        \n_response_1_0_iv_0_0[12]_net_1 , 
        \n_response_1_1_iv_0_0[30]_net_1 , 
        \n_response_1_1_iv_0_0[21]_net_1 , 
        \n_response_1_1_iv_0_0[24]_net_1 , 
        \n_response_1_1_iv_0_0[16]_net_1 , 
        \n_response_1_1_iv_0_0[29]_net_1 , 
        \n_response_1_1_iv_0_0[19]_net_1 , 
        \n_response_1_1_iv_0_0[22]_net_1 , 
        \n_response_1_1_iv_0_0[27]_net_1 , 
        \n_response_1_1_iv_0_0[13]_net_1 , 
        \n_response_123_m_1[1]_net_1 , 
        \n_response_1_1_iv_0_0[34]_net_1 , 
        \state_ns_0_i_o2_0_1_0[0]_net_1 , 
        \state_ns_0_i_o2_0_0[0]_net_1 , 
        n_bus_state_1_sqmuxa_1_i_0_net_1, 
        \n_response_1_1_iv_0_0[14]_net_1 , \state_ns_0_2[3]_net_1 , 
        n_state_2_sqmuxa_0_a6_0_1_net_1, \crc[2] , 
        n_cmd_out_iv_0_o2_2_net_1, \crc[5] , n_cmd_out_iv_0_o2_1, 
        un1_arg_15_5_0, un1_arg_15_4_net_1, 
        \state_ns_i_0_0_0[1]_net_1 , un1_arg_12_9_net_1, 
        n_response_0_sqmuxa_18_0_0_i_1_net_1, 
        n_response_7_sqmuxa_1_0_0_tz_1_net_1, un1_arg_13_i_i_a2_0_13_5, 
        N_3629, n_response_4_sqmuxa, N_285, N_3578, 
        un1_n_bit_0_sqmuxa_i_0, N_1062, N_1061, N_317_1, 
        un1_arg_13_i_i_a2_0_12, N_337, \n_response_123_m[7]_net_1 , 
        \n_response_123_m[3]_net_1 , \n_response_123_m[2]_net_1 , 
        N_3624, N_360, N_631, \n_response_1_0_iv_0_0[5]_net_1 , 
        \n_response_159_m[0] , \n_response_159_m[7]_net_1 , N_89, 
        \n_response_1_0_iv_0_0_2[4]_net_1 , n_state_2_sqmuxa, N_3688_i, 
        \bus_state_ns_0_0_0[2]_net_1 , buffer_under_runlde_0_a6_7, 
        N_4041_i, N_3627, N_3714, N_370, n_response_1_sqmuxa_5, N_2235, 
        N_3685_tz, N_286, \n_response_1_0_iv_0_1[5]_net_1 , 
        \n_response_1_0_iv_2[7]_net_1 , n_cmd_out_iv_0_o2_3_net_1, 
        \n_response_1_0_iv_0_0_4[4]_net_1 , buffer_under_runlde_0_a6_2, 
        buffer_under_runlde_0_a6_8, \state_ns_0_i_o2_0_3[0]_net_1 , 
        \n_response_47_i_2[0]_net_1 , N_140, N_202, un1_arg_12_net_1, 
        un1_arg_15_net_1, \n_response_123_m[0]_net_1 , un86_net_1, 
        N_216, \n_response_1_0_iv_2[3]_net_1 , 
        \n_response_1_0_iv_0_0_3[4]_net_1 , 
        \n_response_1_0_iv_2[6]_net_1 , \n_response_406_m_0[11] , 
        N_3587, N_416, \n_response_392_m[0] , N_3690, 
        \n_response_1_0_iv_0_3[5]_net_1 , N_3707, 
        \n_response_1_0_iv_2[2]_net_1 , N_417, N_145, 
        \n_response_1_0_iv_1[0]_net_1 , 
        \n_response_1_0_iv_0_1[12]_net_1 , N_293, 
        \n_response_360_m[6] , \n_response_49_m[0] , dsd_clkr_net_1, 
        \din[0] , \din[1] , \din[2] , \din[3] , \din[4] , \din[5] , 
        \din[6] , \din[7] , \din[8] , \din[9] , \din[10] , \din[11] , 
        \din[12] , \din[13] , \din[14] , \din[15] , \din[16] , 
        \din[17] , \din[18] , \din[19] , \din[20] , \din[21] , 
        \din[22] , \din[23] , \din[24] , \din[25] , \din[26] , 
        \din[27] , \din[28] , \din[29] , \din[30] , \din[31] , wen, 
        is_last_data, \cnt[5] , \dsd138_ctrl[0] , \dsd138_ctrl[1] , 
        \dsd138_ctrl[2] , i2s_start, master_lrck, spdif_clock_0, 
        dop_clock_0, \source_left[0] , \source_left[1] , 
        \source_left[2] , \source_left[3] , \source_left[4] , 
        \source_left[5] , \source_left[6] , \source_left[7] , 
        \source_left[8] , \source_left[9] , \source_left[10] , 
        \source_left[11] , \source_left[12] , \source_left[13] , 
        \source_left[14] , \source_left[15] , \source_left[16] , 
        \source_left[17] , \source_left[18] , \source_left[19] , 
        \source_left[20] , \source_left[21] , \source_left[22] , 
        \source_left[23] , \source_left[24] , \source_left[25] , 
        \source_left[26] , \source_left[27] , \source_left[28] , 
        \source_left[29] , \source_left[30] , \source_left[31] , 
        \source_right[0] , \source_right[1] , \source_right[2] , 
        \source_right[3] , \source_right[4] , \source_right[5] , 
        \source_right[6] , \source_right[7] , \source_right[8] , 
        \source_right[9] , \source_right[10] , \source_right[11] , 
        \source_right[12] , \source_right[13] , \source_right[14] , 
        \source_right[15] , \source_right[16] , \source_right[17] , 
        \source_right[18] , \source_right[19] , \source_right[20] , 
        \source_right[21] , \source_right[22] , \source_right[23] , 
        \source_right[24] , \source_right[25] , \source_right[26] , 
        \source_right[27] , \source_right[28] , \source_right[29] , 
        \source_right[30] , \source_right[31] , olrck1, olrck2, 
        \dop_right[0] , \dop_right[1] , \dop_right[2] , \dop_right[3] , 
        \dop_right[4] , \dop_right[5] , \dop_right[6] , \dop_right[7] , 
        \dop_right[8] , \dop_right[9] , \dop_right[10] , 
        \dop_right[11] , \dop_right[12] , \dop_right[13] , 
        \dop_right[14] , \dop_right[15] , \dop_left[0] , \dop_left[1] , 
        \dop_left[2] , \dop_left[3] , \dop_left[4] , \dop_left[5] , 
        \dop_left[6] , \dop_left[7] , \dop_left[8] , \dop_left[9] , 
        \dop_left[10] , \dop_left[11] , \dop_left[12] , \dop_left[13] , 
        \dop_left[14] , \dop_left[15] ;
    
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv_1[0]  (.A(
        n_response_0_sqmuxa_1_net_1), .B(\arg[0]_net_1 ), .C(
        \n_response_159_m[0] ), .D(\n_response_392_m[0] ), .Y(
        \n_response_1_0_iv_1[0]_net_1 ));
    CFG3 #( .INIT(8'h0E) )  \n_response_360_1_0[3]  (.A(N_334), .B(
        m42_0_2), .C(\arg[15]_net_1 ), .Y(
        \n_response_360_1_0[3]_net_1 ));
    CFG4 #( .INIT(16'h3100) )  \n_response_123_m_1[1]  (.A(
        n_response_3_sqmuxa_1), .B(\response_i_m[1] ), .C(
        \cccr_func_sel[1]_net_1 ), .D(\state[7]_net_1 ), .Y(
        \n_response_123_m_1[1]_net_1 ));
    SLE response_ret_11 (.D(N_845), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        N_845_reto));
    CFG2 #( .INIT(4'h1) )  \n_response_cnst_4_7_0_.m31_s  (.A(
        \arg[15]_net_1 ), .B(\arg[14]_net_1 ), .Y(m31_s));
    CFG4 #( .INIT(16'hDCEE) )  \n_response_49[2]  (.A(\arg[31]_net_1 ), 
        .B(n_response_49_4_net_1), .C(N_2537), .D(
        \n_response_49_1[2]_net_1 ), .Y(\n_response_49[2]_net_1 ));
    CFG4 #( .INIT(16'h0ACC) )  arg_376 (.A(\arg[30]_net_1 ), .B(
        \arg[31]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_376_net_1));
    SLE \response[39]  (.D(\n_response_1[39] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[39]_net_1 ));
    SLE response_ret_6 (.D(\n_response_cnst_1_m[9] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \n_response_cnst_1_m_reto[9] ));
    CFG2 #( .INIT(4'h8) )  un105_i_a3_0_0 (.A(\arg[31]_net_1 ), .B(
        \state[12]_net_1 ), .Y(N_3641));
    CFG4 #( .INIT(16'hEA00) )  \n_response_123_m[2]  (.A(
        \cccr_func_sel_m[2] ), .B(N_357_i), .C(\response[2]_net_1 ), 
        .D(\state[7]_net_1 ), .Y(\n_response_123_m[2]_net_1 ));
    SLE i_ret_4 (.D(N_3737), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_3737_reto));
    CFG4 #( .INIT(16'h4000) )  un1_arg_12_15_RNI27LT (.A(
        \arg[18]_net_1 ), .B(\arg[14]_net_1 ), .C(\arg[15]_net_1 ), .D(
        N_1062_1_0), .Y(un1_arg_1_1));
    CFG4 #( .INIT(16'h0CAC) )  arg_361 (.A(\arg[15]_net_1 ), .B(
        \arg[16]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_361_net_1));
    CFG4 #( .INIT(16'hF1FD) )  \state_ns_i_0_0_0[1]  (.A(
        \state[1]_net_1 ), .B(\state[0]_net_1 ), .C(N_318), .D(
        n_state13_net_1), .Y(\state_ns_i_0_0_0[1]_net_1 ));
    CFG2 #( .INIT(4'h1) )  n_response_4_sqmuxa_0_a3_0 (.A(
        \arg[11]_net_1 ), .B(\arg[31]_net_1 ), .Y(
        n_response_4_sqmuxa_0_a3_0_net_1));
    CFG3 #( .INIT(8'h01) )  n_response_6_sqmuxa_1 (.A(\arg[13]_net_1 ), 
        .B(\arg[9]_net_1 ), .C(\arg[10]_net_1 ), .Y(
        n_response_6_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'h0020) )  n_state_0_sqmuxa_0_a6_0_a3_1 (.A(
        \ind[2]_net_1 ), .B(\ind[3]_net_1 ), .C(\state[5]_net_1 ), .D(
        \ind[1]_net_1 ), .Y(n_state_0_sqmuxa_0_a6_0_a3_1_net_1));
    CFG4 #( .INIT(16'h88F0) )  \n_response_1_0_iv_1_RNO[0]  (.A(
        \response[0]_net_1 ), .B(\state[8]_net_1 ), .C(
        \n_response_159_m_xx[0]_net_1 ), .D(N_795), .Y(
        \n_response_159_m[0] ));
    CFG4 #( .INIT(16'h009A) )  \n_i_0_iv_0_a6[3]  (.A(\i[3] ), .B(
        \i[2] ), .C(N_276), .D(N_3589_i), .Y(N_3737));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv[8]  (.A(
        \response[8]_net_1 ), .B(\response[7]_net_1 ), .C(N_3595), .D(
        N_845), .Y(\n_response_1[8] ));
    SLE cmden_ret (.D(cmd_out_en_i_reti), .CLK(sdclk_n_1), .EN(
        un96_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        cmd_out_en_i));
    CFG3 #( .INIT(8'h35) )  response_ret_2_RNO_1 (.A(N_4044_i), .B(
        N_66_mux), .C(\arg[15]_net_1 ), .Y(\n_response_360_4_1_1[1] ));
    CFG4 #( .INIT(16'hFFEA) )  \n_response_1_1_iv_0[13]  (.A(
        \n_response_1_1_iv_0_0[13]_net_1 ), .B(\response[12]_net_1 ), 
        .C(N_845), .D(N_145), .Y(\n_response_1[13] ));
    CFG3 #( .INIT(8'h40) )  n_cmd_out29_3 (.A(\i[1] ), .B(\i[0] ), .C(
        N_3736_1), .Y(N_1016_3));
    CFG2 #( .INIT(4'h8) )  un12_n_i_ac0_3 (.A(N_180), .B(\i[2] ), .Y(
        un12_n_i_c3));
    CFG4 #( .INIT(16'hEAAF) )  \state_ns_0_a3_0_a2_i_o3[5]  (.A(
        \ind[3]_net_1 ), .B(N_1386_i), .C(\ind[1]_net_1 ), .D(
        \ind[2]_net_1 ), .Y(N_231));
    CFG4 #( .INIT(16'h0800) )  \n_response_cnst_4_7_0_.m16  (.A(m16_1), 
        .B(N_702_1), .C(\arg[14]_net_1 ), .D(\arg[9]_net_1 ), .Y(
        N_66_mux));
    CFG2 #( .INIT(4'hE) )  \n_response_cnst_4_7_0_.m29_i_o2  (.A(
        \arg[11]_net_1 ), .B(\arg[12]_net_1 ), .Y(N_204));
    CFG4 #( .INIT(16'h7340) )  ind_392 (.A(\state[0]_net_1 ), .B(
        N_3524), .C(\ind[2]_net_1 ), .D(\ind[3]_net_1 ), .Y(
        ind_392_net_1));
    SLE \xo[1]  (.D(\arg[1]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_sound_card_ctrl_1_sqmuxa_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(en49_c));
    CFG4 #( .INIT(16'h0010) )  \state_ns_0_a3_0_a2_4_a3_1[10]  (.A(
        \bus_state[4]_net_1 ), .B(\ind[1]_net_1 ), .C(\ind[0]_net_1 ), 
        .D(\ind[3]_net_1 ), .Y(\state_ns_0_a3_0_a2_4_a3_1[10]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv_0_0_3[4]  (.A(
        \arg[4]_net_1 ), .B(n_response_0_sqmuxa_1_net_1), .C(N_286), 
        .D(N_290), .Y(\n_response_1_0_iv_0_0_3[4]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un1_arg_12 (.A(un1_arg_12_21_net_1), .B(
        un1_arg_12_5_net_1), .C(un1_arg_12_22_net_1), .D(
        un1_arg_12_9_net_1), .Y(un1_arg_12_net_1));
    CFG2 #( .INIT(4'h6) )  \n_i_iv_0_x2[1]  (.A(\i[0] ), .B(\i[1] ), 
        .Y(N_96_i));
    crc7 UCRC (.crc({\crc[6] , \crc[5] , \crc[4] , \crc[3] , \crc[2] , 
        \crc[1] , \crc[0] }), .bit(bit_net_1), .crc_en(crc_en_net_1), 
        .sdclk_n_1(sdclk_n_1), .crc_clr_i(crc_clr_i));
    CFG3 #( .INIT(8'hFE) )  \n_response_1_0_iv[11]  (.A(
        \n_response_cnst_1_m_reto[9] ), .B(\n_response_406_m_reto[11] )
        , .C(\n_response_1_0_iv_0_reto[11] ), .Y(\response[11] ));
    CFG4 #( .INIT(16'h0800) )  n_cmd_out_iv_0_a2 (.A(\state[4]_net_1 ), 
        .B(un1_i_3), .C(N_970), .D(n_cmd_out_iv_0_a2_1_2), .Y(N_147));
    SLE \sound_card_ctrl[5]  (.D(N_3648_i), .CLK(sdclk_n_1), .EN(
        un105_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sound_card_ctrl[5]_net_1 ));
    spdif_tx USPDIF_TX (.source_right({\source_right[31] , 
        \source_right[30] , \source_right[29] , \source_right[28] , 
        \source_right[27] , \source_right[26] , \source_right[25] , 
        \source_right[24] , \source_right[23] , \source_right[22] , 
        \source_right[21] , \source_right[20] , \source_right[19] , 
        \source_right[18] , \source_right[17] , \source_right[16] , 
        \source_right[15] , \source_right[14] , \source_right[13] , 
        \source_right[12] , \source_right[11] , \source_right[10] , 
        \source_right[9] , \source_right[8] }), .source_left({
        \source_left[31] , \source_left[30] , \source_left[29] , 
        \source_left[28] , \source_left[27] , \source_left[26] , 
        \source_left[25] , \source_left[24] , \source_left[23] , 
        \source_left[22] , \source_left[21] , \source_left[20] , 
        \source_left[19] , \source_left[18] , \source_left[17] , 
        \source_left[16] , \source_left[15] , \source_left[14] , 
        \source_left[13] , \source_left[12] , \source_left[11] , 
        \source_left[10] , \source_left[9] , \source_left[8] }), 
        .dop_right({\dop_right[15] , \dop_right[14] , \dop_right[13] , 
        \dop_right[12] , \dop_right[11] , \dop_right[10] , 
        \dop_right[9] , \dop_right[8] , \dop_right[7] , \dop_right[6] , 
        \dop_right[5] , \dop_right[4] , \dop_right[3] , \dop_right[2] , 
        \dop_right[1] , \dop_right[0] }), .dop_left({\dop_left[15] , 
        \dop_left[14] , \dop_left[13] , \dop_left[12] , \dop_left[11] , 
        \dop_left[10] , \dop_left[9] , \dop_left[8] , \dop_left[7] , 
        \dop_left[6] , \dop_left[5] , \dop_left[4] , \dop_left[3] , 
        \dop_left[2] , \dop_left[1] , \dop_left[0] }), .reset_n_i_2(
        reset_n_i_2), .i2s_start(i2s_start), .reset_n_i_0_RNIOUJE(
        reset_n_i_0_RNIOUJE_net_1), .olrck_o(olrck_o), .olrck1(olrck1), 
        .olrck2(olrck2), .use_dsd(use_dsd), .spdif_tx_c(spdif_tx_c), 
        .reset_n_i_i(reset_n_i_i), .spdif_clock_0(spdif_clock_0));
    CFG2 #( .INIT(4'h4) )  \n_response_cnst_4_7_0_.m17_s  (.A(
        \arg[15]_net_1 ), .B(\arg[14]_net_1 ), .Y(m17_s));
    CFG2 #( .INIT(4'h4) )  \n_arg[2]  (.A(\state[0]_net_1 ), .B(
        \arg[1]_net_1 ), .Y(\n_arg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \state_ns_0_i_a2_1[0]  (.A(N_231), .B(
        \state[2]_net_1 ), .Y(N_360));
    CFG4 #( .INIT(16'h0ACC) )  arg_371 (.A(\arg[25]_net_1 ), .B(
        \arg[26]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_371_net_1));
    CFG4 #( .INIT(16'h1020) )  \state_ns_0_a3_2_0[3]  (.A(
        \ind[2]_net_1 ), .B(\ind[3]_net_1 ), .C(\state[5]_net_1 ), .D(
        \ind[1]_net_1 ), .Y(\state_ns_0_a3_2_0_0[3] ));
    CFG4 #( .INIT(16'hCCC8) )  n_state_2_sqmuxa_0_a6_0_1 (.A(N_3692), 
        .B(\state_ns_0_a2_3_1_a6_0_a2_3[0]_net_1 ), .C(\ind[2]_net_1 ), 
        .D(\ind[3]_net_1 ), .Y(n_state_2_sqmuxa_0_a6_0_1_net_1));
    SLE \response[17]  (.D(\n_response_1[17] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[17]_net_1 ));
    SLE \state[6]  (.D(\state_ns[6] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[6]_net_1 ));
    SLE \response[27]  (.D(\n_response_1[27] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[27]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \n_response_cnst_4_7_0_.m42_0_a3_2  (.A(
        N_408), .B(N_10), .C(\arg[11]_net_1 ), .Y(N_336));
    SLE \bus_state[0]  (.D(\bus_state_ns[0] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bus_state[0]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNO[7]  (.A(
        VCC_net_1), .B(\buffer_under_run[7]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[6] ), .S(\buffer_under_run_s[7] ), .Y(), 
        .FCO());
    SLE i_ret_0 (.D(N_3732), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_3732_reto_0));
    CFG4 #( .INIT(16'h1000) )  un1_arg_12_7_0_a2_RNILKEE1 (.A(
        \arg[7]_net_1 ), .B(\arg[4]_net_1 ), .C(un1_arg_0_0), .D(
        un1_arg_12_7), .Y(N_1061));
    CFG1 #( .INIT(2'h1) )  cmden_ret_RNI25J6 (.A(cmd_out_en_i), .Y(
        cmd_out_en_i_i));
    CFG4 #( .INIT(16'h0002) )  n_response_6_sqmuxa (.A(
        n_response_6_sqmuxa_1_net_1), .B(N_4040), .C(\arg[31]_net_1 ), 
        .D(\arg[11]_net_1 ), .Y(n_response_6_sqmuxa_net_1));
    SLE \arg[1]  (.D(\n_arg[1]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[1]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  n_response292 (.A(\arg[9]_net_1 ), .B(
        \arg[13]_net_1 ), .C(N_4040), .D(N_4039), .Y(N_678));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_0_iv_0[7]  (.A(
        \response[6]_net_1 ), .B(\arg[7]_net_1 ), .C(
        n_response_0_sqmuxa_1_net_1), .D(N_845), .Y(
        \n_response_1_0_iv_0[7]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un1_arg_15_RNI324D (.A(un1_arg_12_net_1), 
        .B(un1_arg_15_net_1), .Y(N_3690));
    CFG4 #( .INIT(16'h0A0C) )  \n_response_36[4]  (.A(
        \buffer_under_run[4]_net_1 ), .B(N_1164), .C(N_1166), .D(
        N_1163), .Y(\n_response_36[4]_net_1 ));
    SLE spdif_en (.D(\arg[0]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_spdif_en_1_sqmuxa), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        spdif_en_c));
    CFG2 #( .INIT(4'h4) )  \n_i_0_iv_0_a2_0[5]  (.A(N_3589_i), .B(
        \i[5]_net_1 ), .Y(N_3534));
    CFG4 #( .INIT(16'hFCF8) )  \bus_state_ns_0_0[0]  (.A(N_2266), .B(
        \bus_state[0]_net_1 ), .C(N_3627), .D(N_2265), .Y(
        \bus_state_ns[0] ));
    SLE \arg[17]  (.D(arg_362_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[17]_net_1 ));
    SLE \total_blocks[2]  (.D(\n_total_blocks[2]_net_1 ), .CLK(
        sdclk_n_1), .EN(N_152_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\total_blocks[2]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \i_lm_0[1]  (.A(\n_i_reto[1] ), .B(
        \i_s_reto[1] ), .C(N_3732_reto_2), .Y(\i[1] ));
    CFG3 #( .INIT(8'hBF) )  \state_ns_0_a3_0_a2_i_2[5]  (.A(
        \state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .B(N_4049), .C(
        \ind[0]_net_1 ), .Y(\state_ns_0_a3_0_a2_i_2[5]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  n_state_0_sqmuxa_0_a6_0_a3 (.A(
        \ind[4]_net_1 ), .B(\ind[5]_net_1 ), .C(
        n_state_0_sqmuxa_0_a6_0_a3_1_net_1), .D(\ind[0]_net_1 ), .Y(
        n_state_0_sqmuxa));
    CFG4 #( .INIT(16'h4CCC) )  response_ret_5_RNO_0 (.A(
        n_response_5_sqmuxa_1_1_net_1), .B(\state[10]_net_1 ), .C(
        N_1062), .D(N_1061), .Y(\n_response_406_m_0[11] ));
    SLE in_cmd (.D(\state[1]_net_1 ), .CLK(sdclk_n_1), .EN(
        un97_i_a6_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        in_cmd_net_1));
    SLE \arg[28]  (.D(arg_373_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[28]_net_1 ));
    CFG2 #( .INIT(4'h4) )  un103_i_a2 (.A(N_845), .B(N_181), .Y(N_3762)
        );
    CFG4 #( .INIT(16'h1500) )  \n_response_47_i_a2[0]  (.A(N_4), .B(
        N_1163), .C(\buffer_under_run[0]_net_1 ), .D(N_3592), .Y(
        N_3629));
    CFG3 #( .INIT(8'h10) )  \state_ns_0_a3_0_0[7]  (.A(\arg[21]_net_1 )
        , .B(\arg[17]_net_1 ), .C(N_2175_i_1), .Y(
        \state_ns_0_a3_0_0[7]_net_1 ));
    SLE \arg[26]  (.D(arg_371_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[26]_net_1 ));
    CFG3 #( .INIT(8'hC5) )  \n_response_36[6]  (.A(
        \n_response_36_1_1[6]_net_1 ), .B(\status[6] ), .C(N_1166), .Y(
        \n_response_36[6]_net_1 ));
    CFG4 #( .INIT(16'h45EF) )  \n_response_360_1_0[2]  (.A(
        \arg[14]_net_1 ), .B(\arg[11]_net_1 ), .C(i4_mux_1), .D(N_12), 
        .Y(\n_response_360_1_0[2]_net_1 ));
    SLE \state[2]  (.D(\state_ns[2] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[2]_net_1 ));
    SLE \arg[25]  (.D(arg_370_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[25]_net_1 ));
    CFG2 #( .INIT(4'h8) )  un95_i_a6_0_1 (.A(\i[3] ), .B(\i[2] ), .Y(
        N_3736_1));
    SLE sd_read_start (.D(\state[10]_net_1 ), .CLK(sdclk_n_1), .EN(
        un107_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sd_read_start_net_1));
    SLE response_ret_5 (.D(\n_response_406_m[11] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \n_response_406_m_reto[11] ));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNIP1367[6]  (.A(
        VCC_net_1), .B(\buffer_under_run[6]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[5] ), .S(\buffer_under_run_s[6] ), .Y(), 
        .FCO(\buffer_under_run_cry[6] ));
    CFG4 #( .INIT(16'hBBBA) )  \state_ns_0_4[3]  (.A(
        \state_ns_0_2[3]_net_1 ), .B(N_2181), .C(\state[8]_net_1 ), .D(
        \state[7]_net_1 ), .Y(\state_ns_0_4[3]_net_1 ));
    CFG3 #( .INIT(8'h01) )  bus_state_tr15_6_a2_0 (.A(un1_arg_12_net_1)
        , .B(N_202), .C(un1_arg_15_net_1), .Y(N_1407_i));
    CFG4 #( .INIT(16'hB833) )  \n_response_1_0_iv_0_RNO[5]  (.A(
        N_66_mux), .B(\n_response_1_0_iv_0_m2_6_1[5] ), .C(
        \response[5]_net_1 ), .D(\arg[15]_net_1 ), .Y(N_3572));
    CFG4 #( .INIT(16'h0800) )  n_spdif_en_1_sqmuxa_0_a2 (.A(
        \arg[10]_net_1 ), .B(\arg[11]_net_1 ), .C(N_3592), .D(N_3641), 
        .Y(n_spdif_en_1_sqmuxa));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0[26]  (.A(
        \response[26]_net_1 ), .B(\response[25]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1[26] ));
    CFG4 #( .INIT(16'h0010) )  n_response185 (.A(\arg[10]_net_1 ), .B(
        \arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(\arg[9]_net_1 ), .Y(
        N_1166));
    CFG4 #( .INIT(16'h7350) )  \n_response_1_1_iv_0_0[36]  (.A(
        \response[36]_net_1 ), .B(\response[35]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[36]_net_1 ));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv[35]  (.A(
        \n_response_1_1_iv_0_0[35]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[35] ));
    SLE \buffer_under_run[5]  (.D(\buffer_under_run_s[5] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[5]_net_1 ));
    CFG2 #( .INIT(4'hE) )  n_crc_en_1_sqmuxa_i_o2 (.A(\i[6]_net_1 ), 
        .B(\i[7]_net_1 ), .Y(N_3528));
    SLE i_ret_11 (.D(N_3732), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_3732_reto_2));
    CFG2 #( .INIT(4'h8) )  un12_n_i_ac0_1 (.A(\i[0] ), .B(\i[1] ), .Y(
        N_180));
    SLE \ind[5]  (.D(ind_394_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\ind[5]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \un62_i_a2_0[0]  (.A(\state[3]_net_1 ), .B(
        \state[11]_net_1 ), .C(\state[7]_net_1 ), .Y(N_1697));
    SLE \arg[11]  (.D(arg_356_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[11]_net_1 ));
    CFG4 #( .INIT(16'hEEE2) )  \i_lm_0[2]  (.A(\i_s_reto[2] ), .B(
        N_3732_reto_1), .C(N_74_reto), .D(N_73_reto), .Y(\i[2] ));
    CFG2 #( .INIT(4'h8) )  \state_ns_0_a2_3_1_a6_0_a2[0]  (.A(
        \state_ns_0_a2_3_1_a6_0_a2_3[0]_net_1 ), .B(
        un1_arg_12_22_0_net_1), .Y(N_2222_1_0));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNIN62A4[3]  (.A(
        VCC_net_1), .B(\buffer_under_run[3]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[2] ), .S(\buffer_under_run_s[3] ), .Y(), 
        .FCO(\buffer_under_run_cry[3] ));
    CFG4 #( .INIT(16'h3331) )  \response_RNO[12]  (.A(
        un1_n_bit_0_sqmuxa_i_0), .B(\n_response_1_0_iv_0_1[12]_net_1 ), 
        .C(n_response_1_sqmuxa_net_1), .D(n_state_2_sqmuxa), .Y(
        \n_response_1_0_iv_i[12] ));
    CFG2 #( .INIT(4'h2) )  n_state13 (.A(cmd_q_net_1), .B(cmd_q2_net_1)
        , .Y(n_state13_net_1));
    SLE sd_write_start (.D(N_2938_i), .CLK(sdclk_n_1), .EN(un101_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(sd_write_start_net_1));
    CFG2 #( .INIT(4'h8) )  \n_response_159_m_xx[1]  (.A(
        \n_response_159_m_xx_0[0]_net_1 ), .B(\arg[13]_net_1 ), .Y(
        \n_response_159_m_xx[1]_net_1 ));
    SLE response_ret_2 (.D(\n_response_360[1] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \n_response_360_reto[1] ));
    CFG4 #( .INIT(16'hFEEE) )  \n_response_1_0_iv_0_3[5]  (.A(N_3579), 
        .B(\n_response_1_0_iv_0_1[5]_net_1 ), .C(\state[8]_net_1 ), .D(
        N_3574), .Y(\n_response_1_0_iv_0_3[5]_net_1 ));
    CFG3 #( .INIT(8'hC4) )  n_response_1_sqmuxa (.A(\arg[31]_net_1 ), 
        .B(\state[6]_net_1 ), .C(\arg[28]_net_1 ), .Y(
        n_response_1_sqmuxa_net_1));
    ARI1 #( .INIT(20'h5CCAA) )  \i_cry[0]  (.A(VCC_net_1), .B(\i_0[0] )
        , .C(\i_qxu[0]_net_1 ), .D(GND_net_1), .FCI(i_cry_cy), .S(
        \i_s[0] ), .Y(), .FCO(\i_cry[0]_net_1 ));
    SLE \ind[1]  (.D(ind_390_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\ind[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_arg[6]  (.A(\state[0]_net_1 ), .B(
        \arg[5]_net_1 ), .Y(\n_arg[6]_net_1 ));
    CFG4 #( .INIT(16'hECCC) )  \state_ns_0_i_o2_0_3[0]  (.A(N_317_1), 
        .B(\state_ns_0_i_o2_0_1_0[0]_net_1 ), .C(\ind[3]_net_1 ), .D(
        \state[1]_net_1 ), .Y(\state_ns_0_i_o2_0_3[0]_net_1 ));
    CFG4 #( .INIT(16'hDCEE) )  \n_response_49[3]  (.A(\arg[31]_net_1 ), 
        .B(n_response_49_8_net_1), .C(N_2538), .D(
        \n_response_49_1[3]_net_1 ), .Y(\n_response_49[3]_net_1 ));
    CFG4 #( .INIT(16'h1555) )  n_cmd_out_iv_0_a2_1 (.A(bit_net_1), .B(
        \i[5]_net_1 ), .C(\i[3] ), .D(n_cmd_out_iv_0_a2_7_1_0_net_1), 
        .Y(n_cmd_out_iv_0_a2_1_2));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0080) )  n_state_2_sqmuxa_0_a6_0 (.A(
        \state_ns_0_a3_4_1[3]_net_1 ), .B(un1_arg_12_22_0_net_1), .C(
        n_state_2_sqmuxa_0_a6_0_1_net_1), .D(
        n_state_2_sqmuxa_0_a6_a0_net_1), .Y(n_state_2_sqmuxa));
    CFG4 #( .INIT(16'h0ACC) )  arg_356 (.A(\arg[10]_net_1 ), .B(
        \arg[11]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_356_net_1));
    CFG4 #( .INIT(16'hE3E0) )  \n_response_cnst_4_7_0_.m59  (.A(N_702), 
        .B(\arg[14]_net_1 ), .C(m59_1_1), .D(N_1163), .Y(N_60));
    SLE \buffer_under_run[4]  (.D(\buffer_under_run_s[4] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[4]_net_1 ));
    CFG3 #( .INIT(8'h04) )  no_crc_397_RNO (.A(\state[10]_net_1 ), .B(
        N_1696_i), .C(\state[5]_net_1 ), .Y(N_3747));
    SLE \arg[8]  (.D(\n_arg[8] ), .CLK(sdclk_n_1), .EN(un77), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\arg[8]_net_1 ));
    SLE \cccr_func_sel[2]  (.D(N_3650_i), .CLK(sdclk_n_1), .EN(un87_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cccr_func_sel[2]_net_1 ));
    SLE response_ret_4 (.D(\n_response_1_0_iv_0[11]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\n_response_1_0_iv_0_reto[11] ));
    CFG3 #( .INIT(8'hF1) )  \n_total_blocks[0]  (.A(N_140), .B(
        un1_arg_12_net_1), .C(\arg[0]_net_1 ), .Y(
        \n_total_blocks[0]_net_1 ));
    SLE \response[5]  (.D(\n_response_1[5] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[5]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \state_ns_0_a2_3_10_0_a2[0]  (.A(
        \arg[19]_net_1 ), .B(\arg[27]_net_1 ), .C(\arg[24]_net_1 ), .D(
        \arg[22]_net_1 ), .Y(N_2222_10));
    CFG4 #( .INIT(16'h0CAC) )  arg_362 (.A(\arg[16]_net_1 ), .B(
        \arg[17]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_362_net_1));
    SLE \ind[0]  (.D(ind_389_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\ind[0]_net_1 ));
    CFG4 #( .INIT(16'hFEFA) )  \n_response_1_0_iv_0[5]  (.A(N_3578), 
        .B(\state[9]_net_1 ), .C(\n_response_1_0_iv_0_3[5]_net_1 ), .D(
        N_3572), .Y(\n_response_1[5] ));
    CFG3 #( .INIT(8'hFE) )  n_response_14_sqmuxa_1_o4 (.A(
        \arg[15]_net_1 ), .B(\arg[16]_net_1 ), .C(\arg[14]_net_1 ), .Y(
        N_2721));
    CFG4 #( .INIT(16'hFEEE) )  \n_response_1_1_iv_0[33]  (.A(N_3713), 
        .B(N_3714), .C(\response[33]_net_1 ), .D(N_3595), .Y(
        \n_response_1[33] ));
    CFG4 #( .INIT(16'hFFAE) )  \state_ns_0_i_o2_0_0[0]  (.A(
        \state[11]_net_1 ), .B(\state[0]_net_1 ), .C(n_state13_net_1), 
        .D(N_361), .Y(\state_ns_0_i_o2_0_0[0]_net_1 ));
    CFG3 #( .INIT(8'h08) )  n_state42_0_a2_0_a3 (.A(
        n_state42_0_a2_0_a3_0_net_1), .B(\ind[0]_net_1 ), .C(
        \state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .Y(n_state42));
    SLE response_ret (.D(\n_response_1_0_iv_2[1]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\n_response_1_0_iv_2_reto[1] ));
    SLE \buffer_under_run[2]  (.D(\buffer_under_run_s[2] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[2]_net_1 ));
    CFG4 #( .INIT(16'hFFD0) )  \state_ns_0_i_o2_0_1_0[0]  (.A(
        \ind[0]_net_1 ), .B(\state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .C(
        \state_ns_0_i_a2_0_0[0] ), .D(\state_ns_0_i_o2_0_1[0]_net_1 ), 
        .Y(\state_ns_0_i_o2_0_1_0[0]_net_1 ));
    CFG2 #( .INIT(4'hE) )  n_crc_en_1_sqmuxa_i_o2_RNIT2LH2 (.A(
        n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), .B(un1_i_3), .Y(
        N_213_i));
    CFG4 #( .INIT(16'h4D16) )  \n_response_cnst_4_7_0_.m34  (.A(
        \arg[13]_net_1 ), .B(\arg[9]_net_1 ), .C(\arg[12]_net_1 ), .D(
        \arg[10]_net_1 ), .Y(i4_mux_1));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_0_iv_0[1]  (.A(
        \response[0]_net_1 ), .B(\arg[1]_net_1 ), .C(
        n_response_0_sqmuxa_1_net_1), .D(N_845), .Y(
        \n_response_1_0_iv_0[1]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \i_lm_0[4]  (.A(\i_s[4] ), .B(\n_i[4] ), 
        .C(N_3732), .Y(\i_lm[4] ));
    CFG4 #( .INIT(16'h7FFC) )  n_cmd_out_iv_0_a2_7_1_0 (.A(
        no_crc_net_1), .B(\i[1] ), .C(\i[2] ), .D(\i[0] ), .Y(
        n_cmd_out_iv_0_a2_7_1_0_net_1));
    CFG3 #( .INIT(8'hEC) )  \n_response_1_1_iv_0[14]  (.A(
        \response[13]_net_1 ), .B(\n_response_1_1_iv_0_0[14]_net_1 ), 
        .C(N_845), .Y(\n_response_1[14] ));
    CFG4 #( .INIT(16'h1000) )  \arg_RNI5DQ31[29]  (.A(\arg[29]_net_1 ), 
        .B(\arg[30]_net_1 ), .C(\arg[15]_net_1 ), .D(\arg[14]_net_1 ), 
        .Y(un1_arg_13_i_i_a2_0_13_2));
    ARI1 #( .INIT(20'h45500) )  \state_RNID6CF[12]  (.A(VCC_net_1), .B(
        \state[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(buffer_under_run_cry_cy));
    CLKINT reset_n_i_0_RNIOUJE (.A(reset_n_i_0_0), .Y(
        reset_n_i_0_RNIOUJE_net_1));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_0_iv_0_0[32]  (.A(
        \state[10]_net_1 ), .B(N_3595), .C(\response[32]_net_1 ), .Y(
        \n_response_1_0_iv_0_0[32]_net_1 ));
    CFG4 #( .INIT(16'h00EA) )  n_response_16_sqmuxa_i_0_0 (.A(
        \arg[14]_net_1 ), .B(\arg[12]_net_1 ), .C(\arg[13]_net_1 ), .D(
        N_4054), .Y(n_response_16_sqmuxa_i_0_0_net_1));
    CFG4 #( .INIT(16'hFCFA) )  \n_response_360[7]  (.A(
        \n_response_360_1_0[7]_net_1 ), .B(\response[7]_net_1 ), .C(
        n_response_360_0_net_1), .D(N_709), .Y(
        \n_response_360[7]_net_1 ));
    CFG2 #( .INIT(4'h1) )  un1_arg_12_7_0_a2 (.A(\arg[6]_net_1 ), .B(
        \arg[5]_net_1 ), .Y(un1_arg_12_7));
    CFG3 #( .INIT(8'h80) )  \n_response_cnst_4_7_0_.m42_0_a3_3  (.A(
        N_4), .B(\arg[11]_net_1 ), .C(m42_0_a3_0), .Y(N_337));
    CFG4 #( .INIT(16'hFFEC) )  n_response_0_sqmuxa_18_0_0_i_1 (.A(
        N_685_3), .B(\arg[31]_net_1 ), .C(N_372), .D(N_300), .Y(
        n_response_0_sqmuxa_18_0_0_i_1_net_1));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[21]  (.A(
        \response[21]_net_1 ), .B(\response[20]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[21]_net_1 ));
    CFG4 #( .INIT(16'h880A) )  \n_response_1_0_iv_RNO[0]  (.A(
        \state[12]_net_1 ), .B(\response[0]_net_1 ), .C(N_3587), .D(
        \arg[31]_net_1 ), .Y(\n_response_49_m[0] ));
    CFG4 #( .INIT(16'h00B1) )  \n_response_36[1]  (.A(N_1163), .B(
        n_response_1_sqmuxa_2), .C(\buffer_under_run[1]_net_1 ), .D(
        N_1166), .Y(\n_response_36[1]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  \state_ns_0_a3_0_0_a6_2[8]  (.A(
        \arg[31]_net_1 ), .B(N_2175_i_1), .C(\arg[21]_net_1 ), .D(
        \arg[17]_net_1 ), .Y(\state_ns_0_a3_0_0_a6_2[8]_net_1 ));
    SLE cmd_q (.D(n_cmd_q_net_1), .CLK(sdclk_n_1), .EN(
        un103_i_a6_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        cmd_q_net_1));
    CFG3 #( .INIT(8'hA3) )  \n_response_360[2]  (.A(
        \response[2]_net_1 ), .B(\n_response_360_1_0[2]_net_1 ), .C(
        N_709), .Y(\n_response_360[2]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  \state_ns_0_i_o2_1[0]  (.A(
        \state[2]_net_1 ), .B(N_370), .C(\bus_state[4]_net_1 ), .Y(
        N_216));
    CFG3 #( .INIT(8'h27) )  \n_response_1_0_iv_0_RNO_1[5]  (.A(
        \arg[14]_net_1 ), .B(N_12), .C(N_55), .Y(
        \n_response_1_0_iv_0_m2_6_1_1[5] ));
    CFG4 #( .INIT(16'h0ACC) )  arg_372 (.A(\arg[26]_net_1 ), .B(
        \arg[27]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_372_net_1));
    CFG3 #( .INIT(8'h40) )  \n_response_cnst_4_7_0_.m42_0_a3_0  (.A(
        \arg[13]_net_1 ), .B(N_11), .C(\arg[14]_net_1 ), .Y(N_334));
    CFG3 #( .INIT(8'h28) )  \n_i_0_iv_0_a2_0[2]  (.A(\state[1]_net_1 ), 
        .B(\i[2] ), .C(N_180), .Y(N_74));
    CFG4 #( .INIT(16'h0CAC) )  arg_363 (.A(\arg[17]_net_1 ), .B(
        \arg[18]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_363_net_1));
    CFG2 #( .INIT(4'h8) )  \n_response_159_m_xx_0[0]  (.A(
        \arg[9]_net_1 ), .B(\state[8]_net_1 ), .Y(
        \n_response_159_m_xx_0[0]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \n_response_1_0_iv_0_a3_8[4]  (.A(
        \response[4]_net_1 ), .B(\state[7]_net_1 ), .C(N_357_i), .Y(
        N_290));
    CFG2 #( .INIT(4'h4) )  \n_arg[4]  (.A(\state[0]_net_1 ), .B(
        \arg[3]_net_1 ), .Y(\n_arg[4]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \n_response_1_0_iv_0_a3_7[4]  (.A(
        \state[8]_net_1 ), .B(N_795), .C(\response[4]_net_1 ), .Y(
        N_289));
    CFG2 #( .INIT(4'h2) )  \n_response_360_1_0[7]  (.A(N_60), .B(
        \arg[15]_net_1 ), .Y(\n_response_360_1_0[7]_net_1 ));
    CFG4 #( .INIT(16'h00F8) )  \n_response_1_0_iv_0_0_2[4]  (.A(
        \state[8]_net_1 ), .B(\n_response_cnst_2[6] ), .C(
        \n_response_1_0_iv_0_a3_5_1[4]_net_1 ), .D(N_795), .Y(
        \n_response_1_0_iv_0_0_2[4]_net_1 ));
    SLE \arg[3]  (.D(\n_arg[3]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[3]_net_1 ));
    SLE response_ret_9 (.D(\response[10] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response_reto[10] ));
    SLE \total_blocks[0]  (.D(\n_total_blocks[0]_net_1 ), .CLK(
        sdclk_n_1), .EN(N_152_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\total_blocks[0]_net_1 ));
    CFG4 #( .INIT(16'h7C50) )  \n_i_0_iv_0[4]  (.A(N_3589_i), .B(
        un12_n_i_c4), .C(\i[4]_net_1 ), .D(\state[1]_net_1 ), .Y(
        \n_i[4] ));
    CFG4 #( .INIT(16'h0001) )  \n_response_123_m_RNO[1]  (.A(N_3), .B(
        N_2721), .C(N_243), .D(n_response_0_sqmuxa_18_0_0_i_1_net_1), 
        .Y(N_4041_i));
    CFG2 #( .INIT(4'h1) )  n_response204_1_0_a3_0_a2 (.A(
        \arg[10]_net_1 ), .B(\arg[12]_net_1 ), .Y(N_702_1));
    SLE \arg[10]  (.D(arg_355_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[10]_net_1 ));
    CFG3 #( .INIT(8'h80) )  n_cccr_cd_disable_1_sqmuxa (.A(
        \state[7]_net_1 ), .B(\arg[31]_net_1 ), .C(N_678), .Y(
        n_cccr_cd_disable_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \n_response_1_0_iv[9]  (.A(
        \response_reto[8] ), .B(\n_response_cnst_1_m_reto_1[9] ), .C(
        \n_response_1_0_iv_0_reto[9] ), .D(N_845_reto), .Y(
        \response[9] ));
    CFG4 #( .INIT(16'h3010) )  \i_cry_cy_RNO[0]  (.A(\state[4]_net_1 ), 
        .B(\state[2]_net_1 ), .C(n_state_3_sqmuxa_0_a4_i_c), .D(
        N_213_i), .Y(n_state_3_sqmuxa_0_a4_i_1_0));
    CFG2 #( .INIT(4'h1) )  \n_response_cnst_4_7_0_.m16_1  (.A(
        \arg[11]_net_1 ), .B(\arg[13]_net_1 ), .Y(m16_1));
    CFG2 #( .INIT(4'h4) )  \n_arg[7]  (.A(\state[0]_net_1 ), .B(
        \arg[6]_net_1 ), .Y(\n_arg[7]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \arg_RNI1PTQ[29]  (.A(\arg[30]_net_1 ), .B(
        \arg[29]_net_1 ), .C(\arg[28]_net_1 ), .Y(N_1060));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNIUK1E1[0]  (.A(
        VCC_net_1), .B(\buffer_under_run[0]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        buffer_under_run_cry_cy), .S(\buffer_under_run_s[0] ), .Y(), 
        .FCO(\buffer_under_run_cry[0] ));
    CFG4 #( .INIT(16'h0ACC) )  arg_373 (.A(\arg[27]_net_1 ), .B(
        \arg[28]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_373_net_1));
    SLE \ind[2]  (.D(ind_391_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\ind[2]_net_1 ));
    SLE \ind[3]  (.D(ind_392_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\ind[3]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \bus_state_ns_i_0_a2_0_1[4]  (.A(
        \bus_state[3]_net_1 ), .B(\bus_state[1]_net_1 ), .Y(N_1386_i));
    CFG3 #( .INIT(8'hA3) )  \n_response_cnst_4_7_0_.m48  (.A(N_1163), 
        .B(m48_1_1), .C(\arg[13]_net_1 ), .Y(N_49));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_0_iv_0[6]  (.A(
        \response[5]_net_1 ), .B(\arg[6]_net_1 ), .C(
        n_response_0_sqmuxa_1_net_1), .D(N_845), .Y(
        \n_response_1_0_iv_0[6]_net_1 ));
    CFG2 #( .INIT(4'h1) )  n_cccr_reset_0_sqmuxa_3_0_a2 (.A(
        \arg[9]_net_1 ), .B(\arg[13]_net_1 ), .Y(N_634_1));
    CFG4 #( .INIT(16'h7430) )  ind_390 (.A(\state[0]_net_1 ), .B(
        N_3524), .C(\ind[1]_net_1 ), .D(\ind[0]_net_1 ), .Y(
        ind_390_net_1));
    SLE \response[20]  (.D(\n_response_1[20] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[20]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un102_i_0 (.A(n_sound_card_ctrl_2_sqmuxa), 
        .B(N_355), .Y(un102_i_0_net_1));
    SLE \response[32]  (.D(\n_response_1[32] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[32]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv_2[7]  (.A(
        \state[12]_net_1 ), .B(\n_response_49[7] ), .C(
        \n_response_159_m[7]_net_1 ), .D(
        \n_response_1_0_iv_0[7]_net_1 ), .Y(
        \n_response_1_0_iv_2[7]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_0_iv_0[2]  (.A(
        \response[1] ), .B(\arg[2]_net_1 ), .C(N_845), .D(
        n_response_0_sqmuxa_1_net_1), .Y(
        \n_response_1_0_iv_0[2]_net_1 ));
    CFG2 #( .INIT(4'h2) )  n_response163_2_0_a2 (.A(\arg[9]_net_1 ), 
        .B(\arg[10]_net_1 ), .Y(N_685_3));
    CFG4 #( .INIT(16'h0001) )  un1_state_3_i_a2_0_a6 (.A(
        \state[5]_net_1 ), .B(\state[0]_net_1 ), .C(\state[2]_net_1 ), 
        .D(N_3694), .Y(N_1686_i));
    SLE \response[3]  (.D(\n_response_1[3] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[3]_net_1 ));
    SLE \state[5]  (.D(N_4042_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[5]_net_1 ));
    SLE \sound_card_ctrl[0]  (.D(N_77_i), .CLK(sdclk_n_1), .EN(
        un102_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sound_card_ctrl[0]_net_1 ));
    CFG3 #( .INIT(8'hC4) )  \state_RNIB5A54[4]  (.A(\state[4]_net_1 ), 
        .B(n_state_3_sqmuxa_0_a4_i_0_1), .C(N_213_i), .Y(
        n_state_3_sqmuxa_0_a4_i_0_2));
    CFG3 #( .INIT(8'h01) )  \state_ns_0_a3_3_0_a2[3]  (.A(\i[5]_net_1 )
        , .B(\i[3] ), .C(\i[4]_net_1 ), .Y(N_413));
    CFG4 #( .INIT(16'h8000) )  \state_ns_0_a3_4_1[3]  (.A(
        \state[5]_net_1 ), .B(N_2222_10), .C(\arg[30]_net_1 ), .D(
        \arg[29]_net_1 ), .Y(\state_ns_0_a3_4_1[3]_net_1 ));
    CFG4 #( .INIT(16'hFF40) )  n_cmd_out_iv_0_o2_1_1 (.A(\crc[5] ), .B(
        N_174), .C(N_1013_3), .D(N_163), .Y(n_cmd_out_iv_0_o2_1));
    CFG4 #( .INIT(16'h0F0E) )  n_response_7_sqmuxa_1_0_0 (.A(N_3), .B(
        N_2721), .C(N_678), .D(n_response_7_sqmuxa_1_0_0_tz_1_net_1), 
        .Y(N_795));
    CFG4 #( .INIT(16'h0CAC) )  arg_365 (.A(\arg[19]_net_1 ), .B(
        \arg[20]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_365_net_1));
    CFG3 #( .INIT(8'h01) )  \state_RNO[5]  (.A(N_231), .B(
        \state_ns_0_a3_0_a2_i_2[5]_net_1 ), .C(
        \state_ns_0_a3_0_a2_i_1[5]_net_1 ), .Y(N_4042_i));
    CFG4 #( .INIT(16'hFF10) )  \bus_state_ns_0_0[1]  (.A(N_3666), .B(
        \state[0]_net_1 ), .C(N_3688_i), .D(N_3624), .Y(
        \bus_state_ns[1] ));
    CFG2 #( .INIT(4'h8) )  un1_arg_12_12 (.A(\arg[31]_net_1 ), .B(
        \arg[28]_net_1 ), .Y(un1_arg_12_12_net_1));
    CFG3 #( .INIT(8'hE0) )  \n_total_blocks[2]  (.A(N_140), .B(
        un1_arg_12_net_1), .C(\arg[2]_net_1 ), .Y(
        \n_total_blocks[2]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[19]  (.A(
        \response[19]_net_1 ), .B(\response[18]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[19]_net_1 ));
    SLE \arg[31]  (.D(arg_376_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[31]_net_1 ));
    SLE \ind[4]  (.D(ind_393_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\ind[4]_net_1 ));
    CFG4 #( .INIT(16'hFF08) )  \bus_state_ns_0_0[2]  (.A(
        \state[10]_net_1 ), .B(\bus_state[3]_net_1 ), .C(N_1407_i), .D(
        \bus_state_ns_0_0_0[2]_net_1 ), .Y(\bus_state_ns[2] ));
    CFG3 #( .INIT(8'h01) )  un1_arg_15_0 (.A(\arg[29]_net_1 ), .B(
        \arg[8]_net_1 ), .C(\arg[30]_net_1 ), .Y(un1_arg_15_0_net_1));
    CFG3 #( .INIT(8'h20) )  n_response_360_0 (.A(N_66_mux), .B(N_709), 
        .C(\arg[15]_net_1 ), .Y(n_response_360_0_net_1));
    CFG4 #( .INIT(16'h1F00) )  n_cmd_out4_0_a2_0_a3 (.A(\i[1] ), .B(
        \i[2] ), .C(\i[3] ), .D(n_cmd_out4_0_a2_0_a3_1_net_1), .Y(
        N_970));
    SLE \cccr_func_sel[3]  (.D(N_3649_i), .CLK(sdclk_n_1), .EN(un87_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cccr_func_sel[3]_net_1 ));
    ARI1 #( .INIT(20'h51BE4) )  \i_cry[1]  (.A(N_845_i), .B(
        N_3732_reto_2), .C(\i_s_reto[1] ), .D(\n_i_reto[1] ), .FCI(
        \i_cry[0]_net_1 ), .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0[25]  (.A(
        \response[25]_net_1 ), .B(\response[24]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1[25] ));
    CFG2 #( .INIT(4'h8) )  n_response_14_sqmuxa_1_a4_0_0 (.A(
        \arg[13]_net_1 ), .B(\arg[12]_net_1 ), .Y(N_401));
    CFG4 #( .INIT(16'h60C0) )  \n_i_0_iv_0_a2[5]  (.A(\i[4]_net_1 ), 
        .B(\i[5]_net_1 ), .C(\state[1]_net_1 ), .D(un12_n_i_c4), .Y(
        N_69));
    SLE start_dsd_tx (.D(dop_start), .CLK(dsd_clk_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(start_dsd_tx_net_1));
    CFG3 #( .INIT(8'h16) )  \n_response_cnst_4_7_0_.N_4044_i_1  (.A(
        \arg[12]_net_1 ), .B(\arg[10]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        N_4044_i_1));
    CFG4 #( .INIT(16'h8A80) )  \n_response_1_0_iv_RNO[6]  (.A(
        \state[9]_net_1 ), .B(\response[6]_net_1 ), .C(N_709), .D(
        \n_response_cnst_4[4] ), .Y(\n_response_360_m[6] ));
    CFG4 #( .INIT(16'h4447) )  \n_response_49_1[3]  (.A(
        \response[3]_net_1 ), .B(\arg[31]_net_1 ), .C(N_1166), .D(
        N_706), .Y(\n_response_49_1[3]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  \state_ns_0_a3_3_0_a3_1[3]  (.A(
        \state[9]_net_1 ), .B(\i[1] ), .C(\i[2] ), .D(\i[0] ), .Y(
        \state_ns_0_a3_3_0_a3_1[3]_net_1 ));
    CFG4 #( .INIT(16'h1055) )  sd_write_start_RNO_0 (.A(un101_2_net_1), 
        .B(N_1407_i), .C(\bus_state[3]_net_1 ), .D(\state[10]_net_1 ), 
        .Y(un101_i));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[35]  (.A(
        \response[35]_net_1 ), .B(\response[34]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[35]_net_1 ));
    CFG4 #( .INIT(16'hF5F7) )  \state_ns_0_a3_0_a2_i_1[5]  (.A(
        \state[2]_net_1 ), .B(N_1387_i), .C(\bus_state[4]_net_1 ), .D(
        \ind[2]_net_1 ), .Y(\state_ns_0_a3_0_a2_i_1[5]_net_1 ));
    CFG4 #( .INIT(16'h0CAC) )  arg_375 (.A(\arg[29]_net_1 ), .B(
        \arg[30]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_375_net_1));
    CFG4 #( .INIT(16'h2004) )  \n_response_cnst_4_7_0_.m10  (.A(
        \arg[10]_net_1 ), .B(\arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(
        \arg[9]_net_1 ), .Y(N_11));
    CFG4 #( .INIT(16'h7430) )  ind_393 (.A(\state[0]_net_1 ), .B(
        N_3524), .C(\ind[4]_net_1 ), .D(\ind[3]_net_1 ), .Y(
        ind_393_net_1));
    CFG3 #( .INIT(8'hE0) )  \n_total_blocks[1]  (.A(N_140), .B(
        un1_arg_12_net_1), .C(\arg[1]_net_1 ), .Y(
        \n_total_blocks[1]_net_1 ));
    SLE \xo[0]  (.D(\arg[0]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_sound_card_ctrl_1_sqmuxa_1), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(en45_c));
    CFG2 #( .INIT(4'h8) )  response_ret_10_RNO (.A(N_845), .B(
        \response[9] ), .Y(\response_m_0[9] ));
    SLE \response[35]  (.D(\n_response_1[35] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[35]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \n_response_cnst_4_7_0_.m9_0_a2  (.A(
        \arg[12]_net_1 ), .B(\arg[10]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        N_10));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[27]  (.A(
        \n_response_1_1_iv_0_0[27]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_1_sqmuxa), .Y(\n_response_1[27] ));
    CFG3 #( .INIT(8'h80) )  n_state42_0_a2_0_a3_0 (.A(\ind[1]_net_1 ), 
        .B(\ind[2]_net_1 ), .C(\ind[3]_net_1 ), .Y(
        n_state42_0_a2_0_a3_0_net_1));
    ARI1 #( .INIT(20'h49900) )  \i_s[7]  (.A(VCC_net_1), .B(N_845), .C(
        \i[7]_net_1 ), .D(GND_net_1), .FCI(\i_cry[6]_net_1 ), .S(
        \i_s[7]_net_1 ), .Y(), .FCO());
    CFG3 #( .INIT(8'hE4) )  odata (.A(use_dsd), .B(odata2), .C(odata1), 
        .Y(odata_o));
    CFG4 #( .INIT(16'hAAB8) )  no_crc_397 (.A(no_crc_net_1), .B(N_3747)
        , .C(n_state_0_sqmuxa), .D(N_3707), .Y(no_crc_397_net_1));
    SLE crc_clr (.D(\state[2]_net_1 ), .CLK(sdclk_n_1), .EN(N_144), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(crc_clr_net_1));
    CFG2 #( .INIT(4'h2) )  \n_response_47_i_a2_3[0]  (.A(N_3634_2), .B(
        spdif_en_c), .Y(N_3634));
    CFG4 #( .INIT(16'h0054) )  n_cmd_out_en_iv_0_a6_RNO (.A(N_3528), 
        .B(N_244), .C(n_cmd_out_en_1_sqmuxa_0_0_a3_0_2_1), .D(N_970), 
        .Y(N_967));
    CFG4 #( .INIT(16'hF0F4) )  n_sd_read_start_1_sqmuxa_0_a2_i_o2 (.A(
        \arg[0]_net_1 ), .B(un1_arg_0_1_0_0), .C(\arg[27]_net_1 ), .D(
        \arg[1]_net_1 ), .Y(N_3654));
    CFG3 #( .INIT(8'h04) )  \n_response_1_1_iv_0_a6_1[33]  (.A(
        n_response_1_sqmuxa_net_1), .B(un1_n_bit_0_sqmuxa_i_0), .C(
        \state[0]_net_1 ), .Y(N_3714));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_0_iv_0[3]  (.A(
        \response[2]_net_1 ), .B(\arg[3]_net_1 ), .C(
        n_response_0_sqmuxa_1_net_1), .D(N_845), .Y(
        \n_response_1_0_iv_0[3]_net_1 ));
    CFG4 #( .INIT(16'h0CAC) )  arg_368 (.A(\arg[22]_net_1 ), .B(
        \arg[23]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_368_net_1));
    CLKINT_PRESERVE UCK10 (.A(dsd_clkr_net_1), .Y(dsd_clk_1));
    SLE response_ret_13 (.D(\n_response_cnst_1_m[9] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \n_response_cnst_1_m_reto_1[9] ));
    CFG3 #( .INIT(8'hD0) )  un95_i_0 (.A(\state[4]_net_1 ), .B(N_213_i)
        , .C(N_3685_tz), .Y(un95_i_0_net_1));
    CFG4 #( .INIT(16'h3E0E) )  \n_response_1_0_iv_2_RNO[7]  (.A(
        \sound_card_ctrl[7]_net_1 ), .B(\arg[31]_net_1 ), .C(
        \n_response_49_4_1[7] ), .D(\n_response_49_0[7]_net_1 ), .Y(
        \n_response_49[7] ));
    CFG3 #( .INIT(8'h80) )  \n_response_123_m[6]  (.A(
        \response[6]_net_1 ), .B(\state[7]_net_1 ), .C(N_357_i), .Y(
        \n_response_123_m[6]_net_1 ));
    CFG3 #( .INIT(8'h80) )  n_cmd_out_iv_0_a2_1_1 (.A(N_174), .B(
        \i[2] ), .C(\i[1] ), .Y(n_cmd_out_iv_0_a2_1_1_net_1));
    CFG1 #( .INIT(2'h1) )  crc_clr_RNI9177 (.A(crc_clr_net_1), .Y(
        crc_clr_i));
    CFG4 #( .INIT(16'h0010) )  \un62_i_a2[2]  (.A(\state[7]_net_1 ), 
        .B(\state[6]_net_1 ), .C(N_181), .D(\state[4]_net_1 ), .Y(
        N_1684));
    CFG3 #( .INIT(8'h80) )  \n_response_159_m[3]  (.A(\state[8]_net_1 )
        , .B(N_795), .C(\response[3]_net_1 ), .Y(
        \n_response_159_m[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \n_response_cnst_4_7_0_.m42_0_a3_0_0  (.A(
        \arg[13]_net_1 ), .B(\arg[14]_net_1 ), .Y(m42_0_a3_0));
    CFG2 #( .INIT(4'h4) )  \n_arg[1]  (.A(\state[0]_net_1 ), .B(
        \arg[0]_net_1 ), .Y(\n_arg[1]_net_1 ));
    SLE i_ret_3 (.D(\i_s[0] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_s_reto[0] ));
    CFG3 #( .INIT(8'h80) )  \n_response_1_0_iv_0_a8_3[5]  (.A(
        \response[5]_net_1 ), .B(\state[7]_net_1 ), .C(N_357_i), .Y(
        N_3579));
    CFG3 #( .INIT(8'h20) )  \n_response_123_m_RNO[2]  (.A(
        \cccr_func_sel[2]_net_1 ), .B(\arg[31]_net_1 ), .C(N_612), .Y(
        \cccr_func_sel_m[2] ));
    CFG3 #( .INIT(8'h20) )  n_cmd_out_iv_0_a2_2 (.A(N_1014_3), .B(
        \crc[4] ), .C(N_174), .Y(N_160));
    SLE \response[18]  (.D(\n_response_1[18] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[18]_net_1 ));
    CFG4 #( .INIT(16'h11FC) )  \n_response_1_0_iv_0_RNO_0[5]  (.A(
        \response[5]_net_1 ), .B(\arg[15]_net_1 ), .C(
        \n_response_1_0_iv_0_m2_6_1_1[5] ), .D(N_709), .Y(
        \n_response_1_0_iv_0_m2_6_1[5] ));
    CFG4 #( .INIT(16'hEEEA) )  \n_response_1_1_iv_0[21]  (.A(
        \n_response_1_1_iv_0_0[21]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .D(n_state_1_sqmuxa), .Y(
        \n_response_1[21] ));
    SLE \response[28]  (.D(\n_response_1[28] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[28]_net_1 ));
    CFG3 #( .INIT(8'hDF) )  n_bus_state_1_sqmuxa_1_i_o2_0 (.A(
        \ind[0]_net_1 ), .B(\state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .C(
        \ind[1]_net_1 ), .Y(N_3692));
    CFG4 #( .INIT(16'hCC80) )  \n_response_123_m[0]  (.A(
        n_response_1_sqmuxa_5), .B(\state[7]_net_1 ), .C(
        un1_n_response_3_sqmuxa_i_0), .D(
        \n_response_123_iv_0[0]_net_1 ), .Y(
        \n_response_123_m[0]_net_1 ));
    CFG4 #( .INIT(16'h0CAC) )  arg_364 (.A(\arg[18]_net_1 ), .B(
        \arg[19]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_364_net_1));
    SLE \response[8]  (.D(\n_response_1[8] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[8]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \n_response_123_m_1_RNO[1]  (.A(N_357_i), 
        .B(\response[1] ), .Y(\response_i_m[1] ));
    CFG4 #( .INIT(16'hFFF2) )  \n_response_47_i_2[0]  (.A(N_702), .B(
        en45_c), .C(N_3629), .D(N_3634), .Y(
        \n_response_47_i_2[0]_net_1 ));
    SLE \response[36]  (.D(\n_response_1_1_iv_i[36] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[36]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \n_response_159_m_xx[0]  (.A(
        \n_response_159_m_xx_0[0]_net_1 ), .B(N_204), .C(
        \arg[10]_net_1 ), .Y(\n_response_159_m_xx[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \n_arg_0_a3[8]  (.A(\state[0]_net_1 ), .B(
        \arg[7]_net_1 ), .Y(\n_arg[8] ));
    CFG4 #( .INIT(16'hEA00) )  \n_response_123_m[3]  (.A(
        \cccr_func_sel_m[3] ), .B(N_357_i), .C(\response[3]_net_1 ), 
        .D(\state[7]_net_1 ), .Y(\n_response_123_m[3]_net_1 ));
    CFG4 #( .INIT(16'hB833) )  response_ret_2_RNO (.A(N_4043_i), .B(
        \n_response_360_4_1[1] ), .C(\response[1] ), .D(m31_s), .Y(
        \n_response_360[1] ));
    CFG3 #( .INIT(8'h0D) )  \n_response_cnst_4_7_0_.m54_0_1  (.A(
        \arg[12]_net_1 ), .B(\arg[10]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        m54_0_1));
    CFG2 #( .INIT(4'h4) )  \arg_RNI1JUL[2]  (.A(\state[11]_net_1 ), .B(
        \arg[2]_net_1 ), .Y(N_3650_i));
    CFG4 #( .INIT(16'hFDF7) )  n_state_2_sqmuxa_0_m2 (.A(
        \ind[0]_net_1 ), .B(\ind[1]_net_1 ), .C(
        \state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .D(\ind[2]_net_1 ), .Y(
        N_89));
    CFG3 #( .INIT(8'hCD) )  n_response_0_sqmuxa_18_0_0_i_o2 (.A(
        \arg[13]_net_1 ), .B(N_401), .C(N_204), .Y(N_243));
    CFG3 #( .INIT(8'h14) )  \n_response_cnst_4_7_0_.N_4038_i  (.A(
        \arg[12]_net_1 ), .B(\arg[10]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        N_4038_i));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[29]  (.A(
        \response[29]_net_1 ), .B(\response[28]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[29]_net_1 ));
    CFG3 #( .INIT(8'hE0) )  \n_total_blocks[3]  (.A(N_140), .B(
        un1_arg_12_net_1), .C(\arg[3]_net_1 ), .Y(
        \n_total_blocks[3]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \arg_RNI773M1[11]  (.A(N_4053), .B(
        un1_arg_1_1), .C(\arg[11]_net_1 ), .Y(N_1062));
    CFG4 #( .INIT(16'hEEF0) )  \i_lm_0[5]  (.A(N_69), .B(N_3534), .C(
        \i_s[5] ), .D(N_3732), .Y(\i_lm[5] ));
    CFG4 #( .INIT(16'h0001) )  un1_arg_15_RNO (.A(\arg[4]_net_1 ), .B(
        \arg[5]_net_1 ), .C(\arg[7]_net_1 ), .D(\arg[6]_net_1 ), .Y(
        N_1061_2_0));
    CFG4 #( .INIT(16'h1000) )  \state_RNO[11]  (.A(un1_i_3), .B(
        n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), .C(cccr_reset_net_1), 
        .D(\state[4]_net_1 ), .Y(N_2166_i));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[30]  (.A(
        \n_response_1_1_iv_0_0[30]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_1_sqmuxa), .Y(\n_response_1[30] ));
    CFG4 #( .INIT(16'h8000) )  un1_arg_15_1 (.A(\arg[14]_net_1 ), .B(
        \arg[28]_net_1 ), .C(\arg[31]_net_1 ), .D(\arg[15]_net_1 ), .Y(
        un1_arg_15_1_net_1));
    CFG3 #( .INIT(8'hCA) )  \state_ns_0_a3_0_a2_i_m2[5]  (.A(
        \ind[1]_net_1 ), .B(N_1387_i), .C(N_1386_i), .Y(N_4049));
    CFG2 #( .INIT(4'h7) )  \arg_RNI9BRH[10]  (.A(\arg[11]_net_1 ), .B(
        \arg[10]_net_1 ), .Y(N_4039));
    CFG4 #( .INIT(16'h0001) )  \arg_RNIB02V[8]  (.A(\arg[26]_net_1 ), 
        .B(\arg[8]_net_1 ), .C(\arg[7]_net_1 ), .D(\arg[17]_net_1 ), 
        .Y(un1_arg_13_i_i_a2_0_12_4));
    SLE \arg[12]  (.D(arg_357_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[12]_net_1 ));
    SLE \arg[30]  (.D(arg_375_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[30]_net_1 ));
    SLE \i[5]  (.D(\i_lm[5] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  n_response185_2 (.A(\arg[11]_net_1 ), .B(
        \arg[10]_net_1 ), .Y(N_1166_i_2));
    CFG4 #( .INIT(16'h332E) )  response_ret_2_RNO_0 (.A(
        \n_response_360_4_1_1[1] ), .B(N_709), .C(\response[1] ), .D(
        m31_s), .Y(\n_response_360_4_1[1] ));
    CFG4 #( .INIT(16'hFFC4) )  \n_response_1_0_iv_0_1[12]  (.A(
        \bus_state[3]_net_1 ), .B(\state[10]_net_1 ), .C(N_202), .D(
        \n_response_1_0_iv_0_0[12]_net_1 ), .Y(
        \n_response_1_0_iv_0_1[12]_net_1 ));
    CFG4 #( .INIT(16'h8880) )  \state_ns_0_a3_0[3]  (.A(
        \arg[31]_net_1 ), .B(N_2175_i_1), .C(\arg[21]_net_1 ), .D(
        \arg[17]_net_1 ), .Y(N_2218));
    SLE \buffer_under_run[6]  (.D(\buffer_under_run_s[6] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[6]_net_1 ));
    CFG4 #( .INIT(16'h0CAC) )  arg_374 (.A(\arg[28]_net_1 ), .B(
        \arg[29]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_374_net_1));
    SLE response_ret_1 (.D(\n_response_123_m[1]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\n_response_123_m_reto[1] ));
    SLE \state[4]  (.D(N_2223_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[4]_net_1 ));
    CFG4 #( .INIT(16'h5410) )  \n_response_cnst_4_7_0_.m11_0_a2  (.A(
        \arg[13]_net_1 ), .B(\arg[11]_net_1 ), .C(N_10), .D(N_3), .Y(
        N_12));
    SLE i_ret_12 (.D(\i_s[1] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_s_reto[1] ));
    CFG4 #( .INIT(16'h0001) )  \bus_state_ns_0_0_a2_0[0]  (.A(
        n_state_2_sqmuxa), .B(N_3688_i), .C(\state[0]_net_1 ), .D(
        N_3666), .Y(N_3627));
    CFG3 #( .INIT(8'h04) )  n_state_2_sqmuxa_0_a6_a0_0_0 (.A(
        \ind[1]_net_1 ), .B(\ind[2]_net_1 ), .C(\ind[3]_net_1 ), .Y(
        n_state_2_sqmuxa_0_a6_a0_0));
    CFG4 #( .INIT(16'hFCFA) )  \n_response_360[3]  (.A(
        \n_response_360_1_0[3]_net_1 ), .B(\response[3]_net_1 ), .C(
        n_response_360_0_net_1), .D(N_709), .Y(
        \n_response_360[3]_net_1 ));
    SLE \response[21]  (.D(\n_response_1[21] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[21]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \n_response_1_0_iv_0_a8_2[5]  (.A(
        n_response_6_sqmuxa_net_1), .B(un1_n_response_3_sqmuxa_i_0), 
        .C(\state[7]_net_1 ), .Y(N_3578));
    CFG4 #( .INIT(16'hFFAE) )  n_cmd_q (.A(\state[2]_net_1 ), .B(
        \state[4]_net_1 ), .C(N_213_i), .D(cmd0_net_1), .Y(
        n_cmd_q_net_1));
    CFG4 #( .INIT(16'hF2F0) )  \state_ns_0_2[3]  (.A(N_2186), .B(
        \arg[21]_net_1 ), .C(N_2220), .D(N_2175_i_1), .Y(
        \state_ns_0_2[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  n_sound_card_ctrl_2_sqmuxa_0_a2 (.A(N_706), 
        .B(N_3641), .Y(n_sound_card_ctrl_2_sqmuxa));
    CFG4 #( .INIT(16'h0ACC) )  arg_360 (.A(\arg[14]_net_1 ), .B(
        \arg[15]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_360_net_1));
    CFG4 #( .INIT(16'h6A0E) )  \n_response_cnst_4_7_0_.N_4043_i_1  (.A(
        \arg[10]_net_1 ), .B(\arg[13]_net_1 ), .C(\arg[9]_net_1 ), .D(
        \arg[11]_net_1 ), .Y(N_4043_i_1));
    SLE \response[13]  (.D(\n_response_1[13] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[13]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \bus_state_ns_0_o3[0]  (.A(
        \state[2]_net_1 ), .B(n_state42), .C(\state[0]_net_1 ), .Y(
        N_2266));
    SLE \response[23]  (.D(\n_response_1[23] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[23]_net_1 ));
    CFG3 #( .INIT(8'h53) )  \n_response_36_1_1[6]  (.A(
        \buffer_under_run[6]_net_1 ), .B(N_1164), .C(N_1163), .Y(
        \n_response_36_1_1[6]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  \arg_RNIQJBR2[11]  (.A(
        un1_arg_13_i_i_a2_0_12_4), .B(\arg[11]_net_1 ), .C(N_4053), .D(
        un1_arg_13_i_i_a2_0_12_3), .Y(un1_arg_13_i_i_a2_0_12));
    CFG4 #( .INIT(16'h8000) )  \arg_RNIP4FB6[27]  (.A(
        un1_arg_13_i_i_a2_0_13_4), .B(un1_arg_13_i_i_a2_0_12), .C(
        \arg[27]_net_1 ), .D(un1_arg_13_i_i_a2_0_13_5), .Y(N_140));
    CFG4 #( .INIT(16'h8C80) )  \n_response_1_0_iv_0_a3_4[4]  (.A(
        \response[4]_net_1 ), .B(\state[12]_net_1 ), .C(
        \arg[31]_net_1 ), .D(\n_response_36[4]_net_1 ), .Y(N_286));
    CFG2 #( .INIT(4'h4) )  \state_ns_0_a3_0_a2_4_a2[10]  (.A(N_1387_i), 
        .B(\state[2]_net_1 ), .Y(N_374));
    CFG4 #( .INIT(16'h8000) )  n_sd_read_start_1_sqmuxa_0_a2_i_a2 (.A(
        un1_arg_13_i_i_a2_0_13_4), .B(un1_arg_13_i_i_a2_0_12), .C(
        N_3654), .D(un1_arg_13_i_i_a2_0_13_5), .Y(N_202));
    CFG4 #( .INIT(16'h2230) )  \sound_card_ctrl_RNO[7]  (.A(
        \sound_card_ctrl[7]_net_1 ), .B(\state[11]_net_1 ), .C(
        \arg[7]_net_1 ), .D(n_sound_card_ctrl_2_sqmuxa), .Y(N_3646_i));
    CFG4 #( .INIT(16'h4055) )  sd_read_start_RNO (.A(un107_0_0_net_1), 
        .B(N_202), .C(\bus_state[3]_net_1 ), .D(\state[10]_net_1 ), .Y(
        un107_i));
    CFG4 #( .INIT(16'h8A80) )  \n_response_159_m[7]  (.A(
        \state[8]_net_1 ), .B(\response[7]_net_1 ), .C(N_795), .D(N_3), 
        .Y(\n_response_159_m[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  n_bit_0_sqmuxa (.A(N_213_i), .B(
        \state[4]_net_1 ), .Y(N_845));
    CFG4 #( .INIT(16'h4000) )  n_response_49_4 (.A(\arg[31]_net_1 ), 
        .B(\sound_card_ctrl[2]_net_1 ), .C(N_4), .D(\arg[11]_net_1 ), 
        .Y(n_response_49_4_net_1));
    CFG4 #( .INIT(16'h0A0C) )  \sound_card_ctrl_RNO[6]  (.A(
        \sound_card_ctrl[6]_net_1 ), .B(\arg[6]_net_1 ), .C(
        \state[11]_net_1 ), .D(n_sound_card_ctrl_2_sqmuxa), .Y(
        N_3647_i));
    CFG4 #( .INIT(16'h0100) )  n_response163 (.A(\arg[10]_net_1 ), .B(
        \arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(\arg[9]_net_1 ), .Y(
        N_1164));
    SLE \arg[27]  (.D(arg_372_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[27]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \bus_state_ns_0_o2_i_a2_0_o2[2]  (.A(
        \state[10]_net_1 ), .B(\state[2]_net_1 ), .C(N_1686_i), .D(
        n_state_0_sqmuxa), .Y(N_3666));
    SLE \state[10]  (.D(\state_ns[10] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state[10]_net_1 ));
    CFG4 #( .INIT(16'h5551) )  \response_RNO[37]  (.A(
        \n_response_1_1_iv_0_0[37]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_response_1_sqmuxa_net_1), .D(n_state_0_sqmuxa), .Y(
        \n_response_1_1_iv_i[37] ));
    SLE \sound_card_ctrl[6]  (.D(N_3647_i), .CLK(sdclk_n_1), .EN(
        un105_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sound_card_ctrl[6]_net_1 ));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[28]  (.A(
        \n_response_1_1_iv_0_0[28]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[28] ));
    CFG4 #( .INIT(16'h0015) )  n_crc_en_1_sqmuxa_i_o2_RNIVR871 (.A(
        N_3528), .B(\i[1] ), .C(\i[2] ), .D(\i[3] ), .Y(
        n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1));
    CFG2 #( .INIT(4'h7) )  \arg_RNI0AGF[10]  (.A(\arg[9]_net_1 ), .B(
        \arg[10]_net_1 ), .Y(N_4053));
    CFG2 #( .INIT(4'h2) )  \arg_RNIVGUL[0]  (.A(\arg[0]_net_1 ), .B(
        \state[11]_net_1 ), .Y(N_77_i));
    SLE \state[8]  (.D(\state_ns[8] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[8]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  \state_ns_0_a3_0_a2_4_a3[10]  (.A(
        \state_ns_0_a3_0_a2_4_a3_1[10]_net_1 ), .B(N_374), .C(N_1386_i)
        , .D(N_393), .Y(\state_ns[10] ));
    CFG4 #( .INIT(16'h0CAC) )  arg_370 (.A(\arg[24]_net_1 ), .B(
        \arg[25]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_370_net_1));
    SLE \arg[14]  (.D(arg_359_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[14]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  n_response204_0_a2 (.A(\arg[10]_net_1 ), 
        .B(\arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(\arg[9]_net_1 ), 
        .Y(N_702));
    SLE \arg[5]  (.D(\n_arg[5]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[5]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  un1_state_11_2 (.A(\state[11]_net_1 ), 
        .B(\state[3]_net_1 ), .C(\state[1]_net_1 ), .D(
        \state[2]_net_1 ), .Y(un1_state_11_2_net_1));
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv[1]  (.A(
        \state_reto[9] ), .B(\n_response_360_reto[1] ), .C(
        \n_response_123_m_reto[1] ), .D(\n_response_1_0_iv_2_reto[1] ), 
        .Y(\response[1] ));
    CFG2 #( .INIT(4'hE) )  n_response_14_sqmuxa_1_RNI6I5L (.A(N_659), 
        .B(\arg[31]_net_1 ), .Y(N_357_i));
    CFG3 #( .INIT(8'hAC) )  \n_response_36_0[3]  (.A(
        \buffer_under_run[3]_net_1 ), .B(N_1164), .C(N_1163), .Y(
        N_2538));
    CFG4 #( .INIT(16'h0CAC) )  arg_355 (.A(\arg[9]_net_1 ), .B(
        \arg[10]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_355_net_1));
    CFG4 #( .INIT(16'h0800) )  un1_arg_12_9 (.A(un1_arg_12_12_net_1), 
        .B(un1_arg_12_3_0), .C(N_4053), .D(un1_arg_12_4_net_1), .Y(
        un1_arg_12_9_net_1));
    CFG4 #( .INIT(16'h1D0C) )  \n_response_cnst_4_7_0_.m50_1  (.A(
        \arg[13]_net_1 ), .B(\arg[15]_net_1 ), .C(N_66_mux), .D(N_11), 
        .Y(m50_1_0));
    CFG2 #( .INIT(4'h8) )  sd_write_start_RNO (.A(N_3690), .B(
        \state[10]_net_1 ), .Y(N_2938_i));
    SLE \cccr_func_sel[1]  (.D(N_3651_i), .CLK(sdclk_n_1), .EN(un87_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cccr_func_sel[1]_net_1 ));
    CFG4 #( .INIT(16'h0C04) )  un104_i_a6 (.A(\state[4]_net_1 ), .B(
        un104_i_a6_1_net_1), .C(N_3696), .D(N_213_i), .Y(N_144));
    CFG4 #( .INIT(16'hC0EA) )  \n_response_1_1_iv_0_0[14]  (.A(
        \state[10]_net_1 ), .B(N_3595), .C(\response[14]_net_1 ), .D(
        \bus_state[3]_net_1 ), .Y(\n_response_1_1_iv_0_0[14]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  n_cccr_reset_0_sqmuxa_1_1_i (.A(
        \arg[16]_net_1 ), .B(\arg[14]_net_1 ), .C(\arg[15]_net_1 ), .D(
        \arg[12]_net_1 ), .Y(N_4040));
    CFG3 #( .INIT(8'h60) )  \n_i_0_iv_0_a6_0[3]  (.A(\i[3] ), .B(
        un12_n_i_c3), .C(\state[1]_net_1 ), .Y(N_3738));
    CFG4 #( .INIT(16'h0008) )  \n_response_123_m_RNO[0]  (.A(
        n_response_1_sqmuxa_6_1), .B(N_631), .C(\arg[14]_net_1 ), .D(
        \arg[15]_net_1 ), .Y(n_response_1_sqmuxa_5));
    SLE response_ret_12 (.D(\n_response_1_0_iv_0[9]_net_1 ), .CLK(
        sdclk_n_1), .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\n_response_1_0_iv_0_reto[9] ));
    CFG4 #( .INIT(16'hC080) )  \n_response_1_0_iv_0_0_a3[4]  (.A(
        n_response_4_sqmuxa), .B(un1_n_response_3_sqmuxa_i_0), .C(
        \state[7]_net_1 ), .D(n_response_6_sqmuxa_net_1), .Y(N_285));
    CFG4 #( .INIT(16'hEA00) )  \n_response_123_m[7]  (.A(
        cccr_cd_disable_m), .B(N_357_i), .C(\response[7]_net_1 ), .D(
        \state[7]_net_1 ), .Y(\n_response_123_m[7]_net_1 ));
    SLE \response[34]  (.D(\n_response_1_1_iv_i[34] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[34]_net_1 ));
    SLE \arg[21]  (.D(arg_366_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[21]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un81_i_a2 (.A(\state[2]_net_1 ), .B(
        \state[4]_net_1 ), .Y(N_1699));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[17]  (.A(
        \response[17]_net_1 ), .B(\response[16]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[17]_net_1 ));
    CFG4 #( .INIT(16'h2232) )  \bus_state_ns_0_0[3]  (.A(
        \bus_state_ns_0_a4_1_1[3]_net_1 ), .B(N_2265), .C(
        n_state_2_sqmuxa), .D(N_3688_i), .Y(
        \bus_state_ns_0_0[3]_net_1 ));
    SLE \i[6]  (.D(\i_lm[6] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \n_i_0[6]  (.A(N_3589_i), .B(
        \state[1]_net_1 ), .Y(N_2431));
    CFG4 #( .INIT(16'h0001) )  un1_arg_12_15 (.A(\arg[16]_net_1 ), .B(
        \arg[17]_net_1 ), .C(\arg[13]_net_1 ), .D(\arg[12]_net_1 ), .Y(
        N_1062_1_0));
    CFG4 #( .INIT(16'h0222) )  \state_ns_0_i_a2_2[0]  (.A(
        \state[2]_net_1 ), .B(N_4049), .C(\ind[5]_net_1 ), .D(
        \ind[4]_net_1 ), .Y(N_361));
    SLE \state[1]  (.D(N_2153_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    SLE \arg[19]  (.D(arg_364_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[19]_net_1 ));
    ARI1 #( .INIT(20'h5CCAA) )  \i_cry[2]  (.A(VCC_net_1), .B(\i_0[2] )
        , .C(\i_qxu[2]_net_1 ), .D(GND_net_1), .FCI(\i_cry[1]_net_1 ), 
        .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    CFG3 #( .INIT(8'h1B) )  obck (.A(use_dsd), .B(in_bck_1), .C(
        dsd_clk_1), .Y(obck_o));
    CFG3 #( .INIT(8'h01) )  \n_response_123_m_RNO_0[0]  (.A(
        \arg[31]_net_1 ), .B(\arg[11]_net_1 ), .C(\arg[16]_net_1 ), .Y(
        n_response_1_sqmuxa_6_1));
    SLE \arg[13]  (.D(arg_358_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[13]_net_1 ));
    SLE i_ret (.D(N_2431), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_2431_reto));
    CFG2 #( .INIT(4'h1) )  un83_i_a2 (.A(\state[0]_net_1 ), .B(
        \state[6]_net_1 ), .Y(N_1696_i));
    SLE \response[19]  (.D(\n_response_1[19] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[19]_net_1 ));
    mem_controller uctrl (.din({\din[31] , \din[30] , \din[29] , 
        \din[28] , \din[27] , \din[26] , \din[25] , \din[24] , 
        \din[23] , \din[22] , \din[21] , \din[20] , \din[19] , 
        \din[18] , \din[17] , \din[16] , \din[15] , \din[14] , 
        \din[13] , \din[12] , \din[11] , \din[10] , \din[9] , \din[8] , 
        \din[7] , \din[6] , \din[5] , \din[4] , \din[3] , \din[2] , 
        \din[1] , \din[0] }), .status({\status[7] , \status[6] }), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0({
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0]}), .test_0_HWDATA({
        test_0_HWDATA[31], test_0_HWDATA[30], test_0_HWDATA[29], 
        test_0_HWDATA[28], test_0_HWDATA[27], test_0_HWDATA[26], 
        test_0_HWDATA[25], test_0_HWDATA[24], test_0_HWDATA[23], 
        test_0_HWDATA[22], test_0_HWDATA[21], test_0_HWDATA[20], 
        test_0_HWDATA[19], test_0_HWDATA[18], test_0_HWDATA[17], 
        test_0_HWDATA[16], test_0_HWDATA[15], test_0_HWDATA[14], 
        test_0_HWDATA[13], test_0_HWDATA[12], test_0_HWDATA[11], 
        test_0_HWDATA[10], test_0_HWDATA[9], test_0_HWDATA[8], 
        test_0_HWDATA[7], test_0_HWDATA[6], test_0_HWDATA[5], 
        test_0_HWDATA[4], test_0_HWDATA[3], test_0_HWDATA[2], 
        test_0_HWDATA[1], test_0_HWDATA[0]}), .test_0_HADDR({
        test_0_HADDR[16], test_0_HADDR[15], test_0_HADDR[14], 
        test_0_HADDR[13], test_0_HADDR[12], test_0_HADDR[11], 
        test_0_HADDR[10], test_0_HADDR[9], test_0_HADDR[8], 
        test_0_HADDR[7], test_0_HADDR[6], test_0_HADDR[5], 
        test_0_HADDR[4], test_0_HADDR[3], test_0_HADDR[2]}), 
        .source_right({\source_right[31] , \source_right[30] , 
        \source_right[29] , \source_right[28] , \source_right[27] , 
        \source_right[26] , \source_right[25] , \source_right[24] , 
        \source_right[23] , \source_right[22] , \source_right[21] , 
        \source_right[20] , \source_right[19] , \source_right[18] , 
        \source_right[17] , \source_right[16] , \source_right[15] , 
        \source_right[14] , \source_right[13] , \source_right[12] , 
        \source_right[11] , \source_right[10] , \source_right[9] , 
        \source_right[8] , \source_right[7] , \source_right[6] , 
        \source_right[5] , \source_right[4] , \source_right[3] , 
        \source_right[2] , \source_right[1] , \source_right[0] }), 
        .source_left({\source_left[31] , \source_left[30] , 
        \source_left[29] , \source_left[28] , \source_left[27] , 
        \source_left[26] , \source_left[25] , \source_left[24] , 
        \source_left[23] , \source_left[22] , \source_left[21] , 
        \source_left[20] , \source_left[19] , \source_left[18] , 
        \source_left[17] , \source_left[16] , \source_left[15] , 
        \source_left[14] , \source_left[13] , \source_left[12] , 
        \source_left[11] , \source_left[10] , \source_left[9] , 
        \source_left[8] , \source_left[7] , \source_left[6] , 
        \source_left[5] , \source_left[4] , \source_left[3] , 
        \source_left[2] , \source_left[1] , \source_left[0] }), 
        .dsd138_ctrl({\dsd138_ctrl[2] , \dsd138_ctrl[1] , 
        \dsd138_ctrl[0] }), .test_0_HADDR_i_0(test_0_HADDR_i_0), 
        .test_0_HTRANS_0(test_0_HTRANS_0), .state_0_d0(
        \state[9]_net_1 ), .state_0_0(\state[1]_net_1 ), .bus_state_0(
        \bus_state[3]_net_1 ), .sound_card_ctrl_7(
        \sound_card_ctrl[7]_net_1 ), .sound_card_ctrl_6(
        \sound_card_ctrl[6]_net_1 ), .sound_card_ctrl_5(
        \sound_card_ctrl[5]_net_1 ), .sound_card_ctrl_0(
        \sound_card_ctrl[0]_net_1 ), .sound_card_ctrl_1(
        \sound_card_ctrl[1]_net_1 ), .sound_card_ctrl_2(
        \sound_card_ctrl[2]_net_1 ), .cnt_0(\cnt[5] ), .is_last_data(
        is_last_data), .test_0_HWRITE(test_0_HWRITE), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .wen(wen), 
        .buffer_under_runlde_0_a6_2(buffer_under_runlde_0_a6_2), 
        .sdclk_n_1(sdclk_n_1), .in_bck_1(in_bck_1), .master_lrck(
        master_lrck), .use_dsd(use_dsd), .i2s_start(i2s_start), 
        .mclk_1(mclk_1), .N_4047_i(N_4047_i));
    SLE \response[29]  (.D(\n_response_1[29] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[29]_net_1 ));
    pcm_tx UPCMTX (.source_right({\source_right[31] , 
        \source_right[30] , \source_right[29] , \source_right[28] , 
        \source_right[27] , \source_right[26] , \source_right[25] , 
        \source_right[24] , \source_right[23] , \source_right[22] , 
        \source_right[21] , \source_right[20] , \source_right[19] , 
        \source_right[18] , \source_right[17] , \source_right[16] , 
        \source_right[15] , \source_right[14] , \source_right[13] , 
        \source_right[12] , \source_right[11] , \source_right[10] , 
        \source_right[9] , \source_right[8] , \source_right[7] , 
        \source_right[6] , \source_right[5] , \source_right[4] , 
        \source_right[3] , \source_right[2] , \source_right[1] , 
        \source_right[0] }), .source_left({\source_left[31] , 
        \source_left[30] , \source_left[29] , \source_left[28] , 
        \source_left[27] , \source_left[26] , \source_left[25] , 
        \source_left[24] , \source_left[23] , \source_left[22] , 
        \source_left[21] , \source_left[20] , \source_left[19] , 
        \source_left[18] , \source_left[17] , \source_left[16] , 
        \source_left[15] , \source_left[14] , \source_left[13] , 
        \source_left[12] , \source_left[11] , \source_left[10] , 
        \source_left[9] , \source_left[8] , \source_left[7] , 
        \source_left[6] , \source_left[5] , \source_left[4] , 
        \source_left[3] , \source_left[2] , \source_left[1] , 
        \source_left[0] }), .reset_n_i_1(reset_n_i_1), .start_pcm_tx(
        start_pcm_tx_net_1), .reset_n_i_0_RNIOUJE(
        reset_n_i_0_RNIOUJE_net_1), .olrck2(olrck2), .odata2(odata2), 
        .in_bck_1(in_bck_1), .reset_n_i_i(reset_n_i_i_1));
    dsd_tx UDSDTX (.source_left({\source_left[31] , \source_left[30] , 
        \source_left[29] , \source_left[28] , \source_left[27] , 
        \source_left[26] , \source_left[25] , \source_left[24] , 
        \source_left[23] , \source_left[22] , \source_left[21] , 
        \source_left[20] , \source_left[19] , \source_left[18] , 
        \source_left[17] , \source_left[16] , \source_left[15] , 
        \source_left[14] , \source_left[13] , \source_left[12] , 
        \source_left[11] , \source_left[10] , \source_left[9] , 
        \source_left[8] , \source_left[7] , \source_left[6] , 
        \source_left[5] , \source_left[4] , \source_left[3] , 
        \source_left[2] , \source_left[1] , \source_left[0] }), 
        .source_right({\source_right[31] , \source_right[30] , 
        \source_right[29] , \source_right[28] , \source_right[27] , 
        \source_right[26] , \source_right[25] , \source_right[24] , 
        \source_right[23] , \source_right[22] , \source_right[21] , 
        \source_right[20] , \source_right[19] , \source_right[18] , 
        \source_right[17] , \source_right[16] , \source_right[15] , 
        \source_right[14] , \source_right[13] , \source_right[12] , 
        \source_right[11] , \source_right[10] , \source_right[9] , 
        \source_right[8] , \source_right[7] , \source_right[6] , 
        \source_right[5] , \source_right[4] , \source_right[3] , 
        \source_right[2] , \source_right[1] , \source_right[0] }), 
        .reset_n_i_0(reset_n_i_0), .start_dsd_tx(start_dsd_tx_net_1), 
        .reset_n_i_0_RNIOUJE(reset_n_i_0_RNIOUJE_net_1), .odata1(
        odata1), .olrck1(olrck1), .dsd_clk_1(dsd_clk_1), .reset_n_i_i(
        reset_n_i_i_0));
    CFG3 #( .INIT(8'h35) )  \n_response_49_1_1[6]  (.A(
        \sound_card_ctrl[6]_net_1 ), .B(\response[6]_net_1 ), .C(
        \arg[31]_net_1 ), .Y(\n_response_49_1_1[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[20]  (.A(
        \response[20]_net_1 ), .B(\response[19]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[20]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  n_response155_0_a3 (.A(\arg[10]_net_1 ), 
        .B(\arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(\arg[9]_net_1 ), 
        .Y(N_1163));
    CFG4 #( .INIT(16'h00E4) )  un77_0 (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .C(N_244), .D(N_3538), .Y(un77));
    CFG4 #( .INIT(16'hAAC0) )  \n_response_1_0_iv_0_m2_0[5]  (.A(
        \response[5]_net_1 ), .B(\buffer_under_run[5]_net_1 ), .C(
        N_1163), .D(\arg[31]_net_1 ), .Y(N_3573));
    CFG4 #( .INIT(16'h010F) )  n_bus_state_1_sqmuxa_1_i_0_RNIHI6P (.A(
        \ind[3]_net_1 ), .B(N_89), .C(n_bus_state_1_sqmuxa_1_i_0_net_1)
        , .D(N_2235), .Y(N_3688_i));
    CFG4 #( .INIT(16'hEEE2) )  i_cry_cy_422 (.A(\i_s_reto[2] ), .B(
        N_3732_reto_1), .C(N_74_reto), .D(N_73_reto), .Y(\i_0[2] ));
    CFG4 #( .INIT(16'h0001) )  n_response_0_sqmuxa_1_RNIMG8M (.A(
        \state[10]_net_1 ), .B(n_response_0_sqmuxa_1_net_1), .C(N_3595)
        , .D(N_845), .Y(un1_n_bit_0_sqmuxa_i_0));
    SLE i_ret_2 (.D(\i[0] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_reto[0] ));
    SLE \bus_state[4]  (.D(N_2263_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\bus_state[4]_net_1 ));
    SLE \response[0]  (.D(\n_response_1[0] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[0]_net_1 ));
    CFG3 #( .INIT(8'hDC) )  un75_i (.A(\state[1]_net_1 ), .B(N_3538), 
        .C(\state[0]_net_1 ), .Y(N_3524));
    CFG3 #( .INIT(8'h08) )  n_response_0_sqmuxa_1 (.A(\arg[31]_net_1 ), 
        .B(\state[6]_net_1 ), .C(\arg[28]_net_1 ), .Y(
        n_response_0_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'h1F00) )  \n_response_123_m[1]  (.A(
        n_response_4_sqmuxa), .B(N_4041_i), .C(
        un1_n_response_3_sqmuxa_i_0), .D(\n_response_123_m_1[1]_net_1 )
        , .Y(\n_response_123_m[1]_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  \n_response_47_i[0]  (.A(N_3630), .B(
        \n_response_47_i_2[0]_net_1 ), .C(\sound_card_ctrl[0]_net_1 ), 
        .D(N_706), .Y(N_3587));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[15]  (.A(
        \n_response_1_1_iv_0_0[15]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[15] ));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_1_iv_0_0[13]  (.A(
        \state[10]_net_1 ), .B(N_3595), .C(\response[13]_net_1 ), .D(
        \bus_state[2]_net_1 ), .Y(\n_response_1_1_iv_0_0[13]_net_1 ));
    CFG4 #( .INIT(16'h0C08) )  un1_state_11_1_0_a6 (.A(\ind[3]_net_1 ), 
        .B(\state[5]_net_1 ), .C(N_2235), .D(N_89), .Y(N_3707));
    CFG4 #( .INIT(16'hFF40) )  n_cmd_out_iv_0_o2_2_0 (.A(\crc[2] ), .B(
        N_174), .C(N_1016_3), .D(N_164), .Y(n_cmd_out_iv_0_o2_2_net_1));
    CFG4 #( .INIT(16'h8000) )  un1_arg_15 (.A(N_1061_2_0), .B(
        un1_arg_15_4_net_1), .C(un1_arg_12_22_net_1), .D(
        un1_arg_15_5_0), .Y(un1_arg_15_net_1));
    SLE \sound_card_ctrl[1]  (.D(N_3651_i), .CLK(sdclk_n_1), .EN(
        un102_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sound_card_ctrl[1]_net_1 ));
    CFG4 #( .INIT(16'h0CAC) )  arg_367 (.A(\arg[21]_net_1 ), .B(
        \arg[22]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_367_net_1));
    CFG4 #( .INIT(16'h0ACC) )  arg_358 (.A(\arg[12]_net_1 ), .B(
        \arg[13]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_358_net_1));
    CFG4 #( .INIT(16'hC0EA) )  \state_ns_0[8]  (.A(
        \state_ns_0_a3_0_0_a6_2[8]_net_1 ), .B(N_2181), .C(
        \state[8]_net_1 ), .D(N_2186), .Y(\state_ns[8] ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[31]  (.A(
        \response[31]_net_1 ), .B(\response[30]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[31]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  n_cmd_out_iv_0_a2_5 (.A(N_3736_1), .B(
        N_276), .C(\crc[3] ), .D(N_174), .Y(N_163));
    CFG4 #( .INIT(16'h4C7F) )  \n_response_cnst_4_7_0_.m48_1_1  (.A(
        \arg[9]_net_1 ), .B(\arg[11]_net_1 ), .C(
        n_response_4_sqmuxa_i_1), .D(N_4), .Y(m48_1_1));
    CFG3 #( .INIT(8'hFE) )  \state_ns_0_o3[3]  (.A(\arg[20]_net_1 ), 
        .B(\arg[19]_net_1 ), .C(\arg[18]_net_1 ), .Y(N_2186));
    CFG2 #( .INIT(4'hE) )  \state_ns_0_a2_0_a2_i_o3_0[3]  (.A(
        \ind[4]_net_1 ), .B(\ind[5]_net_1 ), .Y(
        \state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ));
    CFG4 #( .INIT(16'h0111) )  \state_ns_0_1_0[3]  (.A(
        \state[10]_net_1 ), .B(N_2218), .C(
        \state_ns_0_a3_4_1[3]_net_1 ), .D(N_2222_1_0), .Y(
        \state_ns_0_1_0[3]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  n_response_14_sqmuxa_1_tz_1 (.A(
        \arg[16]_net_1 ), .B(\arg[14]_net_1 ), .C(\arg[15]_net_1 ), .D(
        N_401), .Y(n_response_14_sqmuxa_1_tz_1_net_1));
    CFG4 #( .INIT(16'hEEEA) )  \n_response_1_1_iv[22]  (.A(
        \n_response_1_1_iv_0_0[22]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .D(n_state_1_sqmuxa), .Y(
        \n_response_1[22] ));
    CFG4 #( .INIT(16'h0200) )  n_response178 (.A(\arg[10]_net_1 ), .B(
        \arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(\arg[9]_net_1 ), .Y(
        N_1165));
    CFG4 #( .INIT(16'hEEEA) )  \n_response_1_1_iv_0[19]  (.A(
        \n_response_1_1_iv_0_0[19]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .D(n_state_1_sqmuxa), .Y(
        \n_response_1[19] ));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[17]  (.A(
        \n_response_1_1_iv_0_0[17]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[17] ));
    CFG2 #( .INIT(4'h8) )  \state_RNO[12]  (.A(\arg[28]_net_1 ), .B(
        \state[6]_net_1 ), .Y(N_2168_i));
    CFG4 #( .INIT(16'h0ACC) )  arg_354 (.A(\arg[8]_net_1 ), .B(
        \arg[9]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_354_net_1));
    CFG4 #( .INIT(16'h0001) )  \n_response_36_RNO[1]  (.A(N_1166), .B(
        N_1163), .C(N_1165), .D(N_1164), .Y(n_response_1_sqmuxa_2));
    CFG4 #( .INIT(16'h0040) )  n_cmd_out_iv_0_a2_6 (.A(\crc[6] ), .B(
        N_174), .C(\i[3] ), .D(N_3658), .Y(N_164));
    CFG4 #( .INIT(16'h0037) )  cmdo_RNO (.A(n_cmd_out_iv_0_o2_2_net_1), 
        .B(\state[4]_net_1 ), .C(n_cmd_out_iv_0_o2_3_net_1), .D(N_147), 
        .Y(n_cmd_out_iv_i));
    SLE \response[37]  (.D(\n_response_1_1_iv_i[37] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[37]_net_1 ));
    CFG4 #( .INIT(16'hFEFA) )  \n_response_1_0_iv_0[32]  (.A(
        \n_response_1_0_iv_0_0[32]_net_1 ), .B(\response[31]_net_1 ), 
        .C(N_3714), .D(N_845), .Y(\n_response_1[32] ));
    SLE dsd_clkr (.D(dsd_clkr_i_i), .CLK(in_bck_1), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dsd_clkr_net_1));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNI2DD76[5]  (.A(
        VCC_net_1), .B(\buffer_under_run[5]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[4] ), .S(\buffer_under_run_s[5] ), .Y(), 
        .FCO(\buffer_under_run_cry[5] ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[24]  (.A(
        \response[24]_net_1 ), .B(\response[23]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[24]_net_1 ));
    SLE \buffer_under_run[7]  (.D(\buffer_under_run_s[7] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[7]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  n_response_16_sqmuxa_i_0_a3_2 (.A(
        \arg[16]_net_1 ), .B(\arg[15]_net_1 ), .C(N_408), .D(N_229), 
        .Y(N_314));
    CFG3 #( .INIT(8'h20) )  \state_ns_0_a3_2[3]  (.A(\ind[0]_net_1 ), 
        .B(\state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .C(
        \state_ns_0_a3_2_0_0[3] ), .Y(N_2220));
    pcm2dsd DSD138 (.dsd138_ctrl({\dsd138_ctrl[2] , \dsd138_ctrl[1] , 
        \dsd138_ctrl[0] }), .cnt_0(\cnt[5] ), .reset_n_i_i(reset_n_i_i)
        , .in_bck_1(in_bck_1), .use_dsd(use_dsd), .i2s_start(i2s_start)
        , .master_lrck(master_lrck), .spdif_clock_0(spdif_clock_0), 
        .dop_clock_0(dop_clock_0), .start_pcm_tx_2(start_pcm_tx_2), 
        .dop_start(dop_start), .mclk_1(mclk_1));
    SLE i_ret_13 (.D(\n_i[1] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\n_i_reto[1] ));
    CFG4 #( .INIT(16'h30DD) )  \n_response_1_0_iv_2_RNO[1]  (.A(
        \n_response_49_4_1_0[1] ), .B(\arg[31]_net_1 ), .C(
        \n_response_36[1]_net_1 ), .D(\n_response_49_4_1_1[1] ), .Y(
        \n_response_49[1] ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[27]  (.A(
        \response[27]_net_1 ), .B(\response[26]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[27]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  un77_0_a2_0 (.A(\state[1]_net_1 ), .B(
        \i[3] ), .C(\i[4]_net_1 ), .D(\i[5]_net_1 ), .Y(N_3538));
    SLE \bus_state[3]  (.D(\bus_state_ns[3] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bus_state[3]_net_1 ));
    SLE \total_blocks[1]  (.D(\n_total_blocks[1]_net_1 ), .CLK(
        sdclk_n_1), .EN(N_152_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\total_blocks[1]_net_1 ));
    SLE cccr_cd_disable (.D(\arg[7]_net_1 ), .CLK(sdclk_n_1), .EN(
        n_cccr_cd_disable_1_sqmuxa_net_1), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(cccr_cd_disable_net_1));
    CFG3 #( .INIT(8'hA8) )  \state_ns_0_i_a2_0_0_0[0]  (.A(
        \state[2]_net_1 ), .B(N_1387_i), .C(\ind[1]_net_1 ), .Y(
        \state_ns_0_i_a2_0_0[0] ));
    CFG2 #( .INIT(4'h2) )  n_response_3_sqmuxa_1_0_a8_0_a3 (.A(N_612), 
        .B(\arg[31]_net_1 ), .Y(n_response_3_sqmuxa_1));
    CFG4 #( .INIT(16'hFFFE) )  \n_response_1_0_iv[6]  (.A(
        \n_response_360_m[6] ), .B(\n_response_123_m[6]_net_1 ), .C(
        \n_response_1_0_iv_0[6]_net_1 ), .D(
        \n_response_1_0_iv_2[6]_net_1 ), .Y(\n_response_1[6] ));
    CFG4 #( .INIT(16'h1000) )  un1_arg_15_4 (.A(\arg[27]_net_1 ), .B(
        \arg[26]_net_1 ), .C(un1_arg_12_21_net_1), .D(
        un1_arg_15_0_net_1), .Y(un1_arg_15_4_net_1));
    SLE \arg[20]  (.D(arg_365_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[20]_net_1 ));
    CFG4 #( .INIT(16'hFBFA) )  cmd_q2_RNO (.A(\state[2]_net_1 ), .B(
        N_213_i), .C(cmd_q_net_1), .D(\state[4]_net_1 ), .Y(N_341_i));
    CFG2 #( .INIT(4'h4) )  \n_arg[5]  (.A(\state[0]_net_1 ), .B(
        \arg[4]_net_1 ), .Y(\n_arg[5]_net_1 ));
    CFG4 #( .INIT(16'hF888) )  n_response204_0_a2_RNIEUP46 (.A(
        buffer_under_runlde_0_a6_0_1), .B(N_702), .C(N_3690), .D(
        buffer_under_runlde_0_a6_8), .Y(buffer_under_rune));
    CFG4 #( .INIT(16'h88F0) )  \i_lm_0[6]  (.A(N_2431), .B(
        \i[6]_net_1 ), .C(\i_s[6] ), .D(N_3732), .Y(\i_lm[6] ));
    CFG4 #( .INIT(16'h8A80) )  \n_response_1_0_iv_0_a3_11[4]  (.A(
        \state[9]_net_1 ), .B(\response[4]_net_1 ), .C(N_709), .D(
        \n_response_cnst_4[4] ), .Y(N_293));
    CFG3 #( .INIT(8'h20) )  n_cccr_reset_0_sqmuxa_1_0 (.A(
        \arg[31]_net_1 ), .B(N_4039), .C(N_634_1), .Y(
        n_cccr_reset_0_sqmuxa_1_0_net_1));
    CFG3 #( .INIT(8'h08) )  n_state_2_sqmuxa_0_a6_a0 (.A(
        n_state_2_sqmuxa_0_a6_a0_0), .B(\ind[0]_net_1 ), .C(
        \state_ns_0_a2_0_a2_i_o3_0[3]_net_1 ), .Y(
        n_state_2_sqmuxa_0_a6_a0_net_1));
    CFG4 #( .INIT(16'h0222) )  \n_response_cnst_4_7_0_.N_4043_i  (.A(
        N_4043_i_1), .B(N_243), .C(\arg[11]_net_1 ), .D(N_634_1), .Y(
        N_4043_i));
    SLE \i[7]  (.D(\i_lm[7] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    SLE \arg[4]  (.D(\n_arg[4]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  n_response_4_sqmuxa_0_a3_1 (.A(
        \arg[10]_net_1 ), .B(\arg[12]_net_1 ), .Y(
        n_response_4_sqmuxa_i_1));
    SLE \cccr_func_sel[0]  (.D(N_77_i), .CLK(sdclk_n_1), .EN(un87_i), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cccr_func_sel[0]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \n_response_123_m_RNO[3]  (.A(
        \cccr_func_sel[3]_net_1 ), .B(\arg[31]_net_1 ), .C(N_612), .Y(
        \cccr_func_sel_m[3] ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[23]  (.A(
        \response[23]_net_1 ), .B(\response[22]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[23]_net_1 ));
    CFG3 #( .INIT(8'h12) )  \n_i_0_iv_0_a2[2]  (.A(\i[2] ), .B(
        N_3589_i), .C(N_276), .Y(N_73));
    CFG4 #( .INIT(16'h0001) )  un1_arg_15_5_RNO (.A(\arg[3]_net_1 ), 
        .B(\arg[2]_net_1 ), .C(\arg[0]_net_1 ), .D(\arg[1]_net_1 ), .Y(
        N_1061_1_0));
    CFG2 #( .INIT(4'h1) )  n_response_16_sqmuxa_i_0_a2_0 (.A(
        \arg[13]_net_1 ), .B(\arg[14]_net_1 ), .Y(N_408));
    CFG3 #( .INIT(8'h08) )  un96_i_a6_4 (.A(\i[5]_net_1 ), .B(N_3736_1)
        , .C(\i[4]_net_1 ), .Y(N_3736_4));
    SLE \state[0]  (.D(N_154_i), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    SLE \buffer_under_run[0]  (.D(\buffer_under_run_s[0] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  un105_i_a3_0 (.A(\state[12]_net_1 ), .B(
        \state[11]_net_1 ), .Y(N_355));
    CFG4 #( .INIT(16'h8CCC) )  \n_response_1_0_iv_1_RNO_0[0]  (.A(
        \arg[27]_net_1 ), .B(\state[10]_net_1 ), .C(N_1061), .D(N_1062)
        , .Y(\n_response_392_m[0] ));
    CFG4 #( .INIT(16'hC0CA) )  cccr_reset_388 (.A(\arg[3]_net_1 ), .B(
        cccr_reset_net_1), .C(un86_net_1), .D(\state[11]_net_1 ), .Y(
        cccr_reset_388_net_1));
    CFG3 #( .INIT(8'h08) )  \state_ns_0_a3_3_0_a3[3]  (.A(N_413), .B(
        \state_ns_0_a3_3_0_a3_1[3]_net_1 ), .C(N_3528), .Y(N_2221));
    CFG4 #( .INIT(16'h00FE) )  un97_i_a6 (.A(\state[4]_net_1 ), .B(
        \state[0]_net_1 ), .C(\state[1]_net_1 ), .D(N_845), .Y(
        un97_i_a6_net_1));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_0_iv_0[11]  (.A(
        \response[11] ), .B(\response[10] ), .C(N_3595), .D(N_845), .Y(
        \n_response_1_0_iv_0[11]_net_1 ));
    CFG4 #( .INIT(16'h88F0) )  \i_lm_0[7]  (.A(N_2431), .B(
        \i[7]_net_1 ), .C(\i_s[7]_net_1 ), .D(N_3732), .Y(\i_lm[7] ));
    CFG4 #( .INIT(16'hF400) )  \state_RNO[0]  (.A(N_2235), .B(
        \state[5]_net_1 ), .C(N_417), .D(N_416), .Y(N_154_i));
    CFG4 #( .INIT(16'h54BA) )  \n_response_cnst_4_7_0_.m50  (.A(
        \arg[15]_net_1 ), .B(\arg[14]_net_1 ), .C(N_49), .D(m50_1_0), 
        .Y(\n_response_cnst_4[4] ));
    CFG2 #( .INIT(4'hE) )  un1_state_3_i_a2_0_o2_RNI26MI (.A(N_3694), 
        .B(\state[8]_net_1 ), .Y(N_3696));
    CFG3 #( .INIT(8'h01) )  \arg_RNIK9RQ[23]  (.A(\arg[23]_net_1 ), .B(
        \arg[20]_net_1 ), .C(\arg[13]_net_1 ), .Y(
        un1_arg_13_i_i_a2_0_13_1));
    CFG4 #( .INIT(16'h0CAC) )  arg_369 (.A(\arg[23]_net_1 ), .B(
        \arg[24]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_369_net_1));
    CFG4 #( .INIT(16'h0002) )  n_state_1_sqmuxa_0_a6 (.A(
        \state[5]_net_1 ), .B(\ind[2]_net_1 ), .C(\ind[3]_net_1 ), .D(
        N_3692), .Y(n_state_1_sqmuxa));
    CFG2 #( .INIT(4'h8) )  un1_arg_12_22 (.A(N_1062_1_0), .B(
        un1_arg_12_22_0_net_1), .Y(un1_arg_12_22_net_1));
    CFG3 #( .INIT(8'hEC) )  \n_response_1_0_iv_0_1[5]  (.A(
        \response[4]_net_1 ), .B(\n_response_1_0_iv_0_0[5]_net_1 ), .C(
        N_845), .Y(\n_response_1_0_iv_0_1[5]_net_1 ));
    CFG4 #( .INIT(16'h73FF) )  \bus_state_RNO_0[4]  (.A(
        \bus_state[0]_net_1 ), .B(\state[2]_net_1 ), .C(N_1386_i), .D(
        n_state42), .Y(N_2263_i_1));
    CFG3 #( .INIT(8'h75) )  un107_0_0 (.A(N_1684), .B(\state[0]_net_1 )
        , .C(N_979_1), .Y(un107_0_0_net_1));
    CFG4 #( .INIT(16'hFFEC) )  \n_response_1_0_iv[7]  (.A(
        \state[9]_net_1 ), .B(\n_response_123_m[7]_net_1 ), .C(
        \n_response_360[7]_net_1 ), .D(\n_response_1_0_iv_2[7]_net_1 ), 
        .Y(\n_response_1[7] ));
    CFG3 #( .INIT(8'h7F) )  un1_buffer_under_runlto2 (.A(
        \buffer_under_run[2]_net_1 ), .B(\buffer_under_run[1]_net_1 ), 
        .C(\buffer_under_run[0]_net_1 ), .Y(un1_buffer_under_runlt5));
    SLE \state[12]  (.D(N_2168_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[12]_net_1 ));
    SLE \buffer_under_run[3]  (.D(\buffer_under_run_s[3] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[3]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  \arg_RNID8S01[8]  (.A(\arg[0]_net_1 ), 
        .B(un1_arg_0_1_0_0), .C(\arg[8]_net_1 ), .D(\arg[1]_net_1 ), 
        .Y(un1_arg_0_0));
    SLE \bus_state[1]  (.D(\bus_state_ns[1] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bus_state[1]_net_1 ));
    CFG4 #( .INIT(16'hAA4C) )  \n_response_cnst_4_7_0_.m54_0  (.A(
        \arg[11]_net_1 ), .B(m54_0_1), .C(\arg[12]_net_1 ), .D(
        \arg[13]_net_1 ), .Y(m54_0));
    SLE i_ret_8 (.D(N_74), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_74_reto));
    CFG4 #( .INIT(16'h3050) )  n_cmd_out_iv_0_a2_1_0 (.A(\crc[1] ), .B(
        \crc[0] ), .C(\i[3] ), .D(\i[0] ), .Y(
        n_cmd_out_iv_0_a2_1_0_net_1));
    CFG4 #( .INIT(16'hEC00) )  \bus_state_ns_0_0_0[2]  (.A(
        \state[0]_net_1 ), .B(N_3666), .C(data_bus_busy), .D(
        \bus_state[2]_net_1 ), .Y(\bus_state_ns_0_0_0[2]_net_1 ));
    SLE cccr_reset (.D(cccr_reset_388_net_1), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        cccr_reset_net_1));
    CFG2 #( .INIT(4'hE) )  n_cccr_reset_0_sqmuxa_1_1_i_o2 (.A(
        \arg[15]_net_1 ), .B(\arg[16]_net_1 ), .Y(N_4054));
    CFG2 #( .INIT(4'h4) )  \n_arg[3]  (.A(\state[0]_net_1 ), .B(
        \arg[2]_net_1 ), .Y(\n_arg[3]_net_1 ));
    SLE \arg[7]  (.D(\n_arg[7]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[7]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv_2[1]  (.A(
        \state[12]_net_1 ), .B(\n_response_49[1] ), .C(
        \n_response_159_m[1] ), .D(\n_response_1_0_iv_0[1]_net_1 ), .Y(
        \n_response_1_0_iv_2[1]_net_1 ));
    CFG4 #( .INIT(16'h50CC) )  un1_n_response299 (.A(N_3592), .B(N_10), 
        .C(\arg[10]_net_1 ), .D(\arg[13]_net_1 ), .Y(N_631));
    CFG4 #( .INIT(16'hFEFF) )  \state_ns_0[3]  (.A(\state[12]_net_1 ), 
        .B(N_2221), .C(\state_ns_0_4[3]_net_1 ), .D(
        \state_ns_0_1_0[3]_net_1 ), .Y(\state_ns[3] ));
    ARI1 #( .INIT(20'h5CCAA) )  \i_cry[3]  (.A(VCC_net_1), .B(\i_0[3] )
        , .C(\i_qxu[3]_net_1 ), .D(GND_net_1), .FCI(\i_cry[2]_net_1 ), 
        .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    SLE start_pcm_tx (.D(start_pcm_tx_2), .CLK(in_bck_1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(start_pcm_tx_net_1));
    CFG3 #( .INIT(8'hE4) )  \n_response_cnst_4_7_0_.m17_d_d  (.A(
        \arg[15]_net_1 ), .B(N_3), .C(N_66_mux), .Y(m17_d_d));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv[20]  (.A(
        \n_response_1_1_iv_0_0[20]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[20] ));
    SLE \response[2]  (.D(\n_response_1[2] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[2]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \un60_i_a4_0_a2[1]  (.A(
        \bus_state[3]_net_1 ), .B(\bus_state[2]_net_1 ), .Y(N_1387_i));
    CFG4 #( .INIT(16'h0001) )  un1_arg_12_22_0 (.A(\arg[25]_net_1 ), 
        .B(\arg[23]_net_1 ), .C(\arg[20]_net_1 ), .D(\arg[18]_net_1 ), 
        .Y(un1_arg_12_22_0_net_1));
    CFG4 #( .INIT(16'hAA30) )  \n_response_1_0_iv_0_m2_1[5]  (.A(
        \response[5]_net_1 ), .B(\arg[9]_net_1 ), .C(\arg[11]_net_1 ), 
        .D(N_795), .Y(N_3574));
    CFG3 #( .INIT(8'h32) )  n_response_14_sqmuxa_1 (.A(
        n_response_14_sqmuxa_1_tz_1_net_1), .B(N_678), .C(N_3634_2), 
        .Y(N_659));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[16]  (.A(
        \response[16]_net_1 ), .B(\response[15]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[16]_net_1 ));
    SLE cmd0 (.D(cmd_in), .CLK(sdclk_n_i), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(cmd0_net_1));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv[31]  (.A(
        \n_response_1_1_iv_0_0[31]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[31] ));
    CFG4 #( .INIT(16'hFEEE) )  n_cmd_out_iv_0_o2_3 (.A(N_160), .B(
        n_cmd_out_iv_0_o2_1), .C(n_cmd_out_iv_0_a2_1_1_net_1), .D(
        n_cmd_out_iv_0_a2_1_0_net_1), .Y(n_cmd_out_iv_0_o2_3_net_1));
    CFG4 #( .INIT(16'h0123) )  \bus_state_ns_0_1[3]  (.A(
        \state[10]_net_1 ), .B(N_1686_i), .C(N_2266), .D(N_1407_i), .Y(
        \bus_state_ns_0_1[3]_net_1 ));
    ARI1 #( .INIT(20'h5A857) )  \i_cry[6]  (.A(\i[6]_net_1 ), .B(
        \state[4]_net_1 ), .C(n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), 
        .D(un1_i_3), .FCI(\i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(
        \i_cry[6]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_1_iv_0[39]  (.A(
        \response[39]_net_1 ), .B(\response[38]_net_1 ), .C(N_845), .D(
        N_3595), .Y(\n_response_1[39] ));
    CFG4 #( .INIT(16'h7340) )  ind_391 (.A(\state[0]_net_1 ), .B(
        N_3524), .C(\ind[1]_net_1 ), .D(\ind[2]_net_1 ), .Y(
        ind_391_net_1));
    CFG2 #( .INIT(4'h4) )  \cccr_func_sel_RNO[3]  (.A(
        \state[11]_net_1 ), .B(\arg[3]_net_1 ), .Y(N_3649_i));
    CFG3 #( .INIT(8'h80) )  \un62_i_a2_0_RNI0B1C1[0]  (.A(N_1697), .B(
        N_181), .C(N_3589_i), .Y(buffer_under_runlde_0_a6_5));
    CFG4 #( .INIT(16'h4447) )  \n_response_49_1[2]  (.A(
        \response[2]_net_1 ), .B(\arg[31]_net_1 ), .C(N_1166), .D(
        N_706), .Y(\n_response_49_1[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  un95_i_a6_0_1_0_0 (.A(N_3736_4), .B(N_180), 
        .Y(un95_i_a6_0_1_0_0_net_1));
    CFG4 #( .INIT(16'h4505) )  un72_0_a2_RNIJ2U71 (.A(un72), .B(N_612), 
        .C(\state[7]_net_1 ), .D(\arg[31]_net_1 ), .Y(un87_i));
    SLE \response[7]  (.D(\n_response_1[7] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[7]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \arg_RNI0IUL[1]  (.A(\arg[1]_net_1 ), .B(
        \state[11]_net_1 ), .Y(N_3651_i));
    CFG4 #( .INIT(16'hFCAA) )  i_cry_cy_421 (.A(\i_s_reto[3] ), .B(
        N_3738_reto), .C(N_3737_reto), .D(N_3732_reto_0), .Y(\i_0[3] ));
    CFG4 #( .INIT(16'hDDA0) )  \n_response_cnst_4_7_0_.m54_1  (.A(
        \arg[13]_net_1 ), .B(N_4038_i), .C(N_702_1), .D(m54_0), .Y(
        N_55));
    CFG3 #( .INIT(8'h40) )  \n_response_cnst_4_7_0_.m2  (.A(
        \arg[12]_net_1 ), .B(\arg[10]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        N_3));
    SLE \buffer_under_run[1]  (.D(\buffer_under_run_s[1] ), .CLK(
        sdclk_n_1), .EN(buffer_under_rune), .ALn(u8_sb_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\buffer_under_run[1]_net_1 ));
    CFG4 #( .INIT(16'h8F80) )  \n_response_1_0_iv_2_RNO_0[1]  (.A(
        \response[1] ), .B(\state[8]_net_1 ), .C(N_795), .D(
        \n_response_159_m_xx[1]_net_1 ), .Y(\n_response_159_m[1] ));
    CFG4 #( .INIT(16'h0C0D) )  \n_response_1_0_iv_0_0_a3_1[4]  (.A(
        N_612), .B(\arg[31]_net_1 ), .C(N_357_i), .D(N_678), .Y(
        un1_n_response_3_sqmuxa_i_0));
    CFG4 #( .INIT(16'h20A0) )  un103_i_a2_RNIKAPF5 (.A(
        n_state_3_sqmuxa_0_a4_i_0_2), .B(\state[10]_net_1 ), .C(N_3762)
        , .D(N_1407_i), .Y(N_3732));
    CFG2 #( .INIT(4'h8) )  n_sound_card_ctrl_1_sqmuxa_1_0_a2 (.A(N_702)
        , .B(N_3641), .Y(n_sound_card_ctrl_1_sqmuxa_1));
    CFG4 #( .INIT(16'h0CAC) )  arg_357 (.A(\arg[11]_net_1 ), .B(
        \arg[12]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_357_net_1));
    SLE \total_blocks[3]  (.D(\n_total_blocks[3]_net_1 ), .CLK(
        sdclk_n_1), .EN(N_152_i), .ALn(u8_sb_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\total_blocks[3]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \sound_card_ctrl_RNO[5]  (.A(
        \sound_card_ctrl[5]_net_1 ), .B(\arg[3]_net_1 ), .C(
        \state[11]_net_1 ), .D(n_sound_card_ctrl_2_sqmuxa), .Y(
        N_3648_i));
    CFG3 #( .INIT(8'hAC) )  \n_response_159[6]  (.A(
        \response[6]_net_1 ), .B(\n_response_cnst_2[6] ), .C(N_795), 
        .Y(\n_response_159[6]_net_1 ));
    SLE \response[6]  (.D(\n_response_1[6] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[6]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  \arg_RNIAJR31[25]  (.A(\arg[18]_net_1 ), 
        .B(\arg[25]_net_1 ), .C(\arg[31]_net_1 ), .D(\arg[28]_net_1 ), 
        .Y(un1_arg_13_i_i_a2_0_12_3));
    CFG4 #( .INIT(16'hFFFE) )  \n_response_1_0_iv_0_0[4]  (.A(
        \n_response_1_0_iv_0_0_4[4]_net_1 ), .B(N_293), .C(N_285), .D(
        \n_response_1_0_iv_0_0_3[4]_net_1 ), .Y(\n_response_1[4] ));
    SLE \arg[18]  (.D(arg_363_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[18]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8000) )  un83_i_a2_RNIH05O4 (.A(N_1696_i), .B(
        buffer_under_runlde_0_a6_2), .C(N_3696), .D(
        buffer_under_runlde_0_a6_7), .Y(buffer_under_runlde_0_a6_8));
    SLE \arg[16]  (.D(arg_361_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[16]_net_1 ));
    dop_gear UDOP (.dop_right({\dop_right[15] , \dop_right[14] , 
        \dop_right[13] , \dop_right[12] , \dop_right[11] , 
        \dop_right[10] , \dop_right[9] , \dop_right[8] , 
        \dop_right[7] , \dop_right[6] , \dop_right[5] , \dop_right[4] , 
        \dop_right[3] , \dop_right[2] , \dop_right[1] , \dop_right[0] })
        , .dop_left({\dop_left[15] , \dop_left[14] , \dop_left[13] , 
        \dop_left[12] , \dop_left[11] , \dop_left[10] , \dop_left[9] , 
        \dop_left[8] , \dop_left[7] , \dop_left[6] , \dop_left[5] , 
        \dop_left[4] , \dop_left[3] , \dop_left[2] , \dop_left[1] , 
        \dop_left[0] }), .source_right({\source_right[31] , 
        \source_right[30] , \source_right[29] , \source_right[28] , 
        \source_right[27] , \source_right[26] , \source_right[25] , 
        \source_right[24] , \source_right[23] , \source_right[22] , 
        \source_right[21] , \source_right[20] , \source_right[19] , 
        \source_right[18] , \source_right[17] , \source_right[16] , 
        \source_right[15] , \source_right[14] , \source_right[13] , 
        \source_right[12] , \source_right[11] , \source_right[10] , 
        \source_right[9] , \source_right[8] , \source_right[7] , 
        \source_right[6] , \source_right[5] , \source_right[4] , 
        \source_right[3] , \source_right[2] , \source_right[1] , 
        \source_right[0] }), .source_left({\source_left[31] , 
        \source_left[30] , \source_left[29] , \source_left[28] , 
        \source_left[27] , \source_left[26] , \source_left[25] , 
        \source_left[24] , \source_left[23] , \source_left[22] , 
        \source_left[21] , \source_left[20] , \source_left[19] , 
        \source_left[18] , \source_left[17] , \source_left[16] , 
        \source_left[15] , \source_left[14] , \source_left[13] , 
        \source_left[12] , \source_left[11] , \source_left[10] , 
        \source_left[9] , \source_left[8] , \source_left[7] , 
        \source_left[6] , \source_left[5] , \source_left[4] , 
        \source_left[3] , \source_left[2] , \source_left[1] , 
        \source_left[0] }), .reset_n_i_3(reset_n_i_3), 
        .reset_n_i_0_RNIOUJE(reset_n_i_0_RNIOUJE_net_1), .use_dsd(
        use_dsd), .i2s_start(i2s_start), .reset_n_i_i(reset_n_i_i_2), 
        .dop_clock_0(dop_clock_0));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNI3LCB3[2]  (.A(
        VCC_net_1), .B(\buffer_under_run[2]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[1] ), .S(\buffer_under_run_s[2] ), .Y(), 
        .FCO(\buffer_under_run_cry[2] ));
    SLE \arg[15]  (.D(arg_360_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[15]_net_1 ));
    CFG2 #( .INIT(4'h9) )  \i_qxu[2]  (.A(N_845), .B(\i[2] ), .Y(
        \i_qxu[2]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  ind_389 (.A(N_3524), .B(\ind[0]_net_1 ), 
        .C(N_342), .Y(ind_389_net_1));
    CFG4 #( .INIT(16'h2002) )  \n_response_cnst_4_7_0_.m42_0_a3  (.A(
        m42_0_a3_0), .B(N_204), .C(\arg[10]_net_1 ), .D(\arg[9]_net_1 )
        , .Y(N_333));
    CFG4 #( .INIT(16'h0080) )  un1_arg_15_5 (.A(\arg[11]_net_1 ), .B(
        N_1061_1_0), .C(un1_arg_15_1_net_1), .D(N_4053), .Y(
        un1_arg_15_5_0));
    CFG1 #( .INIT(2'h1) )  \i_cry_RNO[1]  (.A(N_845), .Y(N_845_i));
    SLE \arg[22]  (.D(arg_367_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[22]_net_1 ));
    SLE \response[12]  (.D(\n_response_1_0_iv_i[12] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[12]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \n_response_360_1[0]  (.A(
        \n_response_360_0[0]_net_1 ), .B(m17_s), .C(N_12), .Y(
        \n_response_360_1[0]_net_1 ));
    SLE \response[22]  (.D(\n_response_1[22] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[22]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \un62_i_a2_1[2]  (.A(\state[12]_net_1 ), .B(
        \state[5]_net_1 ), .Y(N_181));
    CFG3 #( .INIT(8'h57) )  n_crc_en_1_sqmuxa_i_a2_0_o2 (.A(
        \i[5]_net_1 ), .B(\i[3] ), .C(\i[4]_net_1 ), .Y(N_244));
    CFG3 #( .INIT(8'hFD) )  \state_ns_i_0_o2_0[9]  (.A(\arg[21]_net_1 )
        , .B(\arg[28]_net_1 ), .C(\arg[31]_net_1 ), .Y(N_221));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv[29]  (.A(
        \n_response_1_1_iv_0_0[29]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_1_sqmuxa), .Y(\n_response_1[29] ));
    ARI1 #( .INIT(20'h5A857) )  \i_cry[5]  (.A(\i[5]_net_1 ), .B(
        \state[4]_net_1 ), .C(n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), 
        .D(un1_i_3), .FCI(\i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(
        \i_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h8A80) )  \n_response_159_m[2]  (.A(
        \state[8]_net_1 ), .B(\response[2]_net_1 ), .C(N_795), .D(
        N_1166_i_2), .Y(\n_response_159_m[2]_net_1 ));
    CFG2 #( .INIT(4'h1) )  un103_i_a6_0 (.A(\state[9]_net_1 ), .B(
        \state[6]_net_1 ), .Y(un103_i_a6_0_net_1));
    CFG4 #( .INIT(16'h1000) )  un1_arg_12_21_RNI6JIF1 (.A(
        \arg[12]_net_1 ), .B(\arg[16]_net_1 ), .C(
        un1_arg_13_i_i_a2_0_13_1), .D(un1_arg_12_21_net_1), .Y(
        un1_arg_13_i_i_a2_0_13_5));
    CFG4 #( .INIT(16'h7350) )  \n_response_1_0_iv_0_0[12]  (.A(
        \response[12]_net_1 ), .B(\response[11] ), .C(N_3595), .D(
        N_845), .Y(\n_response_1_0_iv_0_0[12]_net_1 ));
    CFG3 #( .INIT(8'h13) )  \n_response_47_i_a2_0[0]  (.A(
        \buffer_under_run[0]_net_1 ), .B(\arg[11]_net_1 ), .C(N_1163), 
        .Y(N_3630));
    SLE \response[30]  (.D(\n_response_1[30] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[30]_net_1 ));
    CFG4 #( .INIT(16'hFF20) )  \state_ns_0_i_o2_0_5[0]  (.A(
        \state[2]_net_1 ), .B(N_1386_i), .C(\ind[2]_net_1 ), .D(
        \ind[3]_net_1 ), .Y(\state_ns_0_i_o2_0[0]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  n_cmd_out_en_iv_0_a6_RNO_0 (.A(
        \i[4]_net_1 ), .B(\i[1] ), .C(\i[2] ), .D(\i[0] ), .Y(
        n_cmd_out_en_1_sqmuxa_0_0_a3_0_2_1));
    SLE \response[4]  (.D(\n_response_1[4] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[4]_net_1 ));
    SLE i_ret_5 (.D(N_3738), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_3738_reto));
    CFG4 #( .INIT(16'h0054) )  un104_i_a6_1 (.A(\state[12]_net_1 ), .B(
        \state[3]_net_1 ), .C(N_1699), .D(\state[9]_net_1 ), .Y(
        un104_i_a6_1_net_1));
    SLE \state[7]  (.D(\state_ns[7] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[7]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \n_response_47_i_a2_3_2[0]  (.A(
        \arg[10]_net_1 ), .B(\arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(
        \arg[9]_net_1 ), .Y(N_3634_2));
    CFG4 #( .INIT(16'hFDFF) )  un101_2 (.A(N_1696_i), .B(N_1699), .C(
        N_979_1), .D(N_1684), .Y(un101_2_net_1));
    CFG4 #( .INIT(16'hECEE) )  un86 (.A(\state[7]_net_1 ), .B(un72), 
        .C(N_4040), .D(n_cccr_reset_0_sqmuxa_1_0_net_1), .Y(un86_net_1)
        );
    CFG4 #( .INIT(16'h0001) )  un1_arg_12_5 (.A(\arg[30]_net_1 ), .B(
        \arg[8]_net_1 ), .C(\arg[7]_net_1 ), .D(\arg[29]_net_1 ), .Y(
        un1_arg_12_5_net_1));
    CFG4 #( .INIT(16'hEEEA) )  \n_response_1_1_iv[16]  (.A(
        \n_response_1_1_iv_0_0[16]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .D(n_state_1_sqmuxa), .Y(
        \n_response_1[16] ));
    SLE \arg[6]  (.D(\n_arg[6]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_123_iv_0[0]  (.A(
        \cccr_func_sel[0]_net_1 ), .B(\response[0]_net_1 ), .C(
        n_response_3_sqmuxa_1), .D(N_357_i), .Y(
        \n_response_123_iv_0[0]_net_1 ));
    CFG4 #( .INIT(16'h0042) )  \n_response_cnst_4_7_0_.N_4044_i  (.A(
        \arg[11]_net_1 ), .B(N_4044_i_1), .C(\arg[12]_net_1 ), .D(
        \arg[13]_net_1 ), .Y(N_4044_i));
    CFG3 #( .INIT(8'h41) )  n_response_0_sqmuxa_18_0_0_i_a3 (.A(
        \arg[11]_net_1 ), .B(\arg[13]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        N_300));
    CFG4 #( .INIT(16'hFFEC) )  \n_response_1_0_iv[3]  (.A(
        \state[9]_net_1 ), .B(\n_response_123_m[3]_net_1 ), .C(
        \n_response_360[3]_net_1 ), .D(\n_response_1_0_iv_2[3]_net_1 ), 
        .Y(\n_response_1[3] ));
    CFG4 #( .INIT(16'h4000) )  \state_ns_i_0_0_a3_0[1]  (.A(
        \state[0]_net_1 ), .B(\i[1] ), .C(\i[2] ), .D(N_318_4), .Y(
        N_318));
    CFG4 #( .INIT(16'h0001) )  n_cmd_out4_0_a2_0_a3_1 (.A(\i[5]_net_1 )
        , .B(\i[4]_net_1 ), .C(N_3528), .D(crc_en_net_1), .Y(
        n_cmd_out4_0_a2_0_a3_1_net_1));
    CFG1 #( .INIT(2'h1) )  reset_n_i_0_RNIOUJE_0 (.A(
        reset_n_i_0_RNIOUJE_net_1), .Y(N_4047_i));
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv_2[2]  (.A(
        \state[12]_net_1 ), .B(\n_response_49[2]_net_1 ), .C(
        \n_response_159_m[2]_net_1 ), .D(
        \n_response_1_0_iv_0[2]_net_1 ), .Y(
        \n_response_1_0_iv_2[2]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[18]  (.A(
        \response[18]_net_1 ), .B(\response[17]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[18]_net_1 ));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[23]  (.A(
        \n_response_1_1_iv_0_0[23]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[23] ));
    CFG3 #( .INIT(8'h14) )  \n_response_cnst_4_7_0_.m17_d_s  (.A(
        \arg[15]_net_1 ), .B(\arg[13]_net_1 ), .C(\arg[11]_net_1 ), .Y(
        m17_d_s));
    SLE \arg[9]  (.D(arg_354_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[9]_net_1 ));
    SLE \sound_card_ctrl[2]  (.D(N_3650_i), .CLK(sdclk_n_1), .EN(
        un102_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sound_card_ctrl[2]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  un1_buffer_under_runlto5 (.A(
        \buffer_under_run[3]_net_1 ), .B(un1_buffer_under_runlt5), .C(
        \buffer_under_run[5]_net_1 ), .D(\buffer_under_run[4]_net_1 ), 
        .Y(un1_buffer_under_runlt7));
    CFG4 #( .INIT(16'hFEFC) )  \n_response_1_1_iv[10]  (.A(
        \response_reto[10] ), .B(\response_m_0_reto[9] ), .C(
        \n_response_cnst_1_m_reto_0[9] ), .D(N_3595_reto), .Y(
        \response[10] ));
    ARI1 #( .INIT(20'h4BF3F) )  \i_cry_cy[0]  (.A(\state[10]_net_1 ), 
        .B(N_1407_i), .C(N_3762), .D(n_state_3_sqmuxa_0_a4_i_1_0), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(i_cry_cy));
    CFG4 #( .INIT(16'hFFCE) )  cmden_ret_RNO (.A(\state[4]_net_1 ), .B(
        \state[0]_net_1 ), .C(N_213_i), .D(N_3724), .Y(
        cmd_out_en_i_reti));
    CFG4 #( .INIT(16'h0010) )  n_response_16_sqmuxa_i_0_a3_1_RNIDVSG (
        .A(N_314), .B(n_response_16_sqmuxa_i_0_0_net_1), .C(N_659), .D(
        N_313), .Y(N_709));
    CFG3 #( .INIT(8'h20) )  \n_response_123_m_RNO[7]  (.A(
        cccr_cd_disable_net_1), .B(\arg[31]_net_1 ), .C(N_678), .Y(
        cccr_cd_disable_m));
    SLE \state[11]  (.D(N_2166_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[11]_net_1 ));
    SLE \response[15]  (.D(\n_response_1[15] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[15]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \n_response_1_1_iv_0_o2[14]  (.A(
        \state[8]_net_1 ), .B(\state[7]_net_1 ), .C(\state[12]_net_1 ), 
        .D(\state[9]_net_1 ), .Y(N_3595));
    CFG4 #( .INIT(16'hFFEA) )  \n_response_1_0_iv_0_0_4[4]  (.A(
        \n_response_1_0_iv_0_0_2[4]_net_1 ), .B(N_845), .C(
        \response[3]_net_1 ), .D(N_289), .Y(
        \n_response_1_0_iv_0_0_4[4]_net_1 ));
    SLE \response[25]  (.D(\n_response_1[25] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[25]_net_1 ));
    CFG3 #( .INIT(8'h04) )  \n_response_cnst_4_7_0_.m3_0_a2  (.A(
        \arg[12]_net_1 ), .B(\arg[10]_net_1 ), .C(\arg[9]_net_1 ), .Y(
        N_4));
    CFG4 #( .INIT(16'h0100) )  \state_ns_0_i_a2_6[0]  (.A(un1_i_3), .B(
        n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), .C(cccr_reset_net_1), 
        .D(\state[4]_net_1 ), .Y(N_370));
    CFG4 #( .INIT(16'h8000) )  \state_ns_0_i_a3_0_0[0]  (.A(
        \arg[30]_net_1 ), .B(\arg[29]_net_1 ), .C(N_2222_10), .D(
        N_2222_1_0), .Y(N_2235));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[22]  (.A(
        \response[22]_net_1 ), .B(\response[21]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[22]_net_1 ));
    SLE \arg[24]  (.D(arg_369_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[24]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0[38]  (.A(
        \response[38]_net_1 ), .B(\response[37]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1[38] ));
    CFG3 #( .INIT(8'hFB) )  n_cmd_out_iv_0_o2_2 (.A(\i[2] ), .B(\i[0] )
        , .C(\i[1] ), .Y(N_3658));
    CFG4 #( .INIT(16'hFFAE) )  \state_ns_0_i_o2_1_0[0]  (.A(
        \state[11]_net_1 ), .B(\state[0]_net_1 ), .C(n_state13_net_1), 
        .D(N_374), .Y(\state_ns_0_i_o2_1[0]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \state_ns_0_a3_0_a2_4_a2_0[10]  (.A(
        \ind[5]_net_1 ), .B(\ind[4]_net_1 ), .C(\ind[2]_net_1 ), .Y(
        N_393));
    CFG2 #( .INIT(4'h9) )  \i_qxu[3]  (.A(N_845), .B(\i[3] ), .Y(
        \i_qxu[3]_net_1 ));
    CFG2 #( .INIT(4'h1) )  un72_0_a2 (.A(\state[7]_net_1 ), .B(
        \state[11]_net_1 ), .Y(un72));
    CFG4 #( .INIT(16'h0CAC) )  arg_359 (.A(\arg[13]_net_1 ), .B(
        \arg[14]_net_1 ), .C(un77), .D(\state[0]_net_1 ), .Y(
        arg_359_net_1));
    CFG2 #( .INIT(4'h1) )  \arg_RNIBS4D[2]  (.A(\arg[3]_net_1 ), .B(
        \arg[2]_net_1 ), .Y(un1_arg_0_1_0_0));
    CFG4 #( .INIT(16'hAF8C) )  \bus_state_RNO[4]  (.A(
        \bus_state[4]_net_1 ), .B(\state[0]_net_1 ), .C(N_2263_i_1), 
        .D(N_3666), .Y(N_2263_i));
    CFG4 #( .INIT(16'hAAD8) )  \n_response_49_0[7]  (.A(N_1166), .B(
        \status[7] ), .C(N_2541), .D(N_702), .Y(
        \n_response_49_0[7]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \n_response_1_0_iv_0_a3_5_1[4]  (.A(
        \state[8]_net_1 ), .B(\arg[12]_net_1 ), .C(N_4053), .Y(
        \n_response_1_0_iv_0_a3_5_1[4]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \i_lm_0_RNIJLDN[0]  (.A(\i[0] ), .B(\i[1] ), 
        .Y(N_276));
    CFG4 #( .INIT(16'h4000) )  un1_arg_12_4 (.A(\arg[26]_net_1 ), .B(
        \arg[14]_net_1 ), .C(\arg[15]_net_1 ), .D(\arg[11]_net_1 ), .Y(
        un1_arg_12_4_net_1));
    SLE i_ret_6 (.D(\i_s[3] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_s_reto[3] ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[30]  (.A(
        \response[30]_net_1 ), .B(\response[29]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[30]_net_1 ));
    SLE i_ret_1 (.D(N_3732), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_3732_reto));
    CFG4 #( .INIT(16'h0111) )  \i_RNIU6CA1[6]  (.A(\i[6]_net_1 ), .B(
        \i[7]_net_1 ), .C(\i[5]_net_1 ), .D(\i[4]_net_1 ), .Y(un1_i_3));
    CFG4 #( .INIT(16'h0001) )  un1_arg_12_21 (.A(\arg[22]_net_1 ), .B(
        \arg[24]_net_1 ), .C(\arg[21]_net_1 ), .D(\arg[19]_net_1 ), .Y(
        un1_arg_12_21_net_1));
    CFG2 #( .INIT(4'h7) )  reset_n_i_0_inst_1 (.A(
        \sound_card_ctrl[7]_net_1 ), .B(u8_sb_0_HPMS_READY), .Y(
        reset_n_i_0_0));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv[18]  (.A(
        \n_response_1_1_iv_0_0[18]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_0_sqmuxa), .Y(\n_response_1[18] ));
    SLE \arg[29]  (.D(arg_374_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[29]_net_1 ));
    SLE response_ret_7 (.D(N_3595), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        N_3595_reto));
    CFG3 #( .INIT(8'h45) )  \n_response_cnst_4_7_0_.m59_1_1  (.A(
        \arg[13]_net_1 ), .B(N_11), .C(\arg[14]_net_1 ), .Y(m59_1_1));
    SLE \arg[23]  (.D(arg_368_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[23]_net_1 ));
    CFG4 #( .INIT(16'hD050) )  \state_ns_0_i_o2_0_1[0]  (.A(
        \ind[2]_net_1 ), .B(\ind[0]_net_1 ), .C(N_374), .D(N_1386_i), 
        .Y(\state_ns_0_i_o2_0_1[0]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un1_state_3_i_a2_0_o2 (.A(\state[10]_net_1 )
        , .B(\state[11]_net_1 ), .Y(N_3694));
    sd_data UD100 (.total_blocks({\total_blocks[3]_net_1 , 
        \total_blocks[2]_net_1 , \total_blocks[1]_net_1 , 
        \total_blocks[0]_net_1 }), .sd_data_out({sd_data_out[3], 
        sd_data_out[2], sd_data_out[1], sd_data_out[0]}), .din({
        \din[31] , \din[30] , \din[29] , \din[28] , \din[27] , 
        \din[26] , \din[25] , \din[24] , \din[23] , \din[22] , 
        \din[21] , \din[20] , \din[19] , \din[18] , \din[17] , 
        \din[16] , \din[15] , \din[14] , \din[13] , \din[12] , 
        \din[11] , \din[10] , \din[9] , \din[8] , \din[7] , \din[6] , 
        \din[5] , \din[4] , \din[3] , \din[2] , \din[1] , \din[0] }), 
        .sd_data_in({sd_data_in[3], sd_data_in[2], sd_data_in[1], 
        sd_data_in[0]}), .status_0(\status[7] ), .in_cmd(in_cmd_net_1), 
        .sd_read_start(sd_read_start_net_1), .sd_write_start(
        sd_write_start_net_1), .data_bus_busy(data_bus_busy), .wen(wen)
        , .is_last_data(is_last_data), .sdclk_n_1(sdclk_n_1), 
        .sdclk_n_i(sdclk_n_i), .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY), 
        .data_out_en_ret_fast_i(data_out_en_ret_fast_i), 
        .sd_data_out_en_i_i(sd_data_out_en_i_i));
    CFG4 #( .INIT(16'hC0EA) )  \state_ns_0[7]  (.A(
        \state_ns_0_a3_0_0[7]_net_1 ), .B(N_2181), .C(\state[7]_net_1 )
        , .D(N_2186), .Y(\state_ns[7] ));
    CFG4 #( .INIT(16'h4000) )  n_response_49_8 (.A(\arg[31]_net_1 ), 
        .B(\sound_card_ctrl[5]_net_1 ), .C(N_4), .D(\arg[11]_net_1 ), 
        .Y(n_response_49_8_net_1));
    CFG3 #( .INIT(8'h40) )  \state_ns_i_0_0_a3_1[1]  (.A(N_413), .B(
        N_244), .C(N_393), .Y(N_317_1));
    SLE \response[16]  (.D(\n_response_1[16] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[16]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  n_response_4_sqmuxa_0_a3 (.A(
        n_response_4_sqmuxa_0_a3_0_net_1), .B(n_response_4_sqmuxa_i_1), 
        .C(N_634_1), .D(N_2721), .Y(n_response_4_sqmuxa));
    CFG3 #( .INIT(8'h47) )  \n_response_1_0_iv_2_RNO_0[7]  (.A(
        \response[7]_net_1 ), .B(\arg[31]_net_1 ), .C(N_702), .Y(
        \n_response_49_4_1[7] ));
    SLE \response[26]  (.D(\n_response_1[26] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[26]_net_1 ));
    CFG3 #( .INIT(8'h04) )  \n_response_cnst_2_0_a2_0_0_a2[4]  (.A(
        \arg[9]_net_1 ), .B(\arg[11]_net_1 ), .C(\arg[10]_net_1 ), .Y(
        \n_response_cnst_2[6] ));
    CFG3 #( .INIT(8'h20) )  bus_state_tr15_6_a2_0_RNIDF5E1 (.A(
        \state[10]_net_1 ), .B(N_1407_i), .C(\bus_state[3]_net_1 ), .Y(
        N_152_i));
    CFG2 #( .INIT(4'hB) )  n_bus_state_1_sqmuxa_1_i_0 (.A(
        n_state_0_sqmuxa), .B(\state[5]_net_1 ), .Y(
        n_bus_state_1_sqmuxa_1_i_0_net_1));
    CFG4 #( .INIT(16'h0080) )  n_cmd_out19_3 (.A(\i[3] ), .B(\i[0] ), 
        .C(\i[1] ), .D(\i[2] ), .Y(N_1014_3));
    SLE \response[38]  (.D(\n_response_1[38] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[38]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \n_response_cnst_4_7_0_.m29_i_a2  (.A(
        \arg[11]_net_1 ), .B(\arg[12]_net_1 ), .Y(N_372));
    CFG4 #( .INIT(16'hFCAA) )  \i_lm_0[3]  (.A(\i_s_reto[3] ), .B(
        N_3738_reto), .C(N_3737_reto), .D(N_3732_reto_0), .Y(\i[3] ));
    CFG2 #( .INIT(4'h2) )  \un62_i_a2_0_RNIOB2U[0]  (.A(N_1697), .B(
        \state[10]_net_1 ), .Y(N_979_1));
    CFG2 #( .INIT(4'h8) )  n_state_2_sqmuxa_0_a6_0_RNIOENU (.A(
        un1_n_bit_0_sqmuxa_i_0), .B(n_state_2_sqmuxa), .Y(
        \n_response_cnst_1_m[9] ));
    CFG4 #( .INIT(16'h8000) )  \state_ns_0_a3_0_a2_0_a3[2]  (.A(
        \state[1]_net_1 ), .B(\i[1] ), .C(\i[2] ), .D(N_318_4), .Y(
        \state_ns[2] ));
    CFG4 #( .INIT(16'hEAC0) )  \n_response_1_0_iv_2[6]  (.A(
        \state[8]_net_1 ), .B(\state[12]_net_1 ), .C(
        \n_response_49[6]_net_1 ), .D(\n_response_159[6]_net_1 ), .Y(
        \n_response_1_0_iv_2[6]_net_1 ));
    CFG4 #( .INIT(16'hE000) )  un96_i_a6 (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(N_180), .D(N_3736_4), .Y(N_3745));
    SLE response_ret_10 (.D(\response_m_0[9] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response_m_0_reto[9] ));
    CFG2 #( .INIT(4'h4) )  \state_RNIDPNF[6]  (.A(\arg[28]_net_1 ), .B(
        \state[6]_net_1 ), .Y(N_2175_i_1));
    CFG2 #( .INIT(4'h1) )  \state_RNI3NHD[8]  (.A(\state[7]_net_1 ), 
        .B(\state[8]_net_1 ), .Y(N_3589_i));
    CFG4 #( .INIT(16'h0020) )  n_response221_0_a2_0_a2 (.A(
        \arg[10]_net_1 ), .B(\arg[12]_net_1 ), .C(\arg[11]_net_1 ), .D(
        \arg[9]_net_1 ), .Y(N_706));
    CFG4 #( .INIT(16'h0501) )  un1_state_11_2_RNIDT123 (.A(
        un1_state_11_2_net_1), .B(\state[4]_net_1 ), .C(N_3707), .D(
        N_213_i), .Y(un1_state_11_i));
    CFG4 #( .INIT(16'hFEF0) )  un105_i_0 (.A(N_706), .B(N_702), .C(
        N_355), .D(N_3641), .Y(un105_i_0_net_1));
    SLE \sound_card_ctrl[7]  (.D(N_3646_i), .CLK(sdclk_n_1), .EN(
        un105_i_0_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sound_card_ctrl[7]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[15]  (.A(
        \response[15]_net_1 ), .B(\response[14]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[15]_net_1 ));
    SLE bit (.D(\response[39]_net_1 ), .CLK(sdclk_n_1), .EN(N_845), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(bit_net_1));
    CFG3 #( .INIT(8'h08) )  n_cmd_out_en_iv_0_a6 (.A(\state[4]_net_1 ), 
        .B(N_967), .C(crc_en_net_1), .Y(N_3724));
    CFG3 #( .INIT(8'h10) )  \state_RNIGASC1[9]  (.A(\state[9]_net_1 ), 
        .B(\state[2]_net_1 ), .C(n_state_3_sqmuxa_0_a4_i_c), .Y(
        n_state_3_sqmuxa_0_a4_i_0_1));
    ARI1 #( .INIT(20'h5A857) )  \i_cry[4]  (.A(\i[4]_net_1 ), .B(
        \state[4]_net_1 ), .C(n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), 
        .D(un1_i_3), .FCI(\i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(
        \i_cry[4]_net_1 ));
    SLE \arg[0]  (.D(N_342), .CLK(sdclk_n_1), .EN(un77), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\arg[0]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  n_response338_0_a3 (.A(\arg[13]_net_1 ), 
        .B(N_685_3), .C(N_2721), .D(N_372), .Y(N_612));
    SLE i_ret_10 (.D(\i_s[2] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_s_reto[2] ));
    CFG4 #( .INIT(16'h0020) )  n_cmd_out14_3 (.A(\i[3] ), .B(\i[0] ), 
        .C(\i[1] ), .D(\i[2] ), .Y(N_1013_3));
    SLE \bus_state[2]  (.D(\bus_state_ns[2] ), .CLK(sdclk_n_1), .EN(
        VCC_net_1), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bus_state[2]_net_1 ));
    CFG4 #( .INIT(16'h1115) )  \response_RNO[34]  (.A(
        \n_response_1_1_iv_0_0[34]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(\state[0]_net_1 ), .D(n_state_1_sqmuxa), .Y(
        \n_response_1_1_iv_i[34] ));
    CFG2 #( .INIT(4'hD) )  \bus_state_RNIHNAV[3]  (.A(
        \state[10]_net_1 ), .B(\bus_state[3]_net_1 ), .Y(
        n_state_3_sqmuxa_0_a4_i_c));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_1_iv_0_0[28]  (.A(
        \response[28]_net_1 ), .B(\response[27]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[28]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \n_response_1_0_iv_0_0[5]  (.A(
        \state[12]_net_1 ), .B(\arg[5]_net_1 ), .C(N_3573), .D(
        n_response_0_sqmuxa_1_net_1), .Y(
        \n_response_1_0_iv_0_0[5]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \n_response_36_0[2]  (.A(
        \buffer_under_run[2]_net_1 ), .B(N_1165), .C(N_1163), .Y(
        N_2537));
    SLE i_ret_9 (.D(N_3732), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_3732_reto_1));
    SLE cmdo (.D(n_cmd_out_iv_i), .CLK(sdclk_n_1), .EN(un95_i_0_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(cmd_out));
    SLE \state[3]  (.D(\state_ns[3] ), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[3]_net_1 ));
    SLE cmd_q2 (.D(N_341_i), .CLK(sdclk_n_1), .EN(un103_i_a6_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(cmd_q2_net_1));
    CFG4 #( .INIT(16'hF0EE) )  un95_i_0_tz (.A(\state[0]_net_1 ), .B(
        \state[4]_net_1 ), .C(un95_i_a6_0_1_0_0_net_1), .D(
        \state[1]_net_1 ), .Y(N_3685_tz));
    CFG3 #( .INIT(8'h80) )  \n_response_1_1_iv_0_a2[13]  (.A(
        \state[10]_net_1 ), .B(N_202), .C(\bus_state[3]_net_1 ), .Y(
        N_145));
    SLE i_ret_7 (.D(N_73), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(N_73_reto));
    CFG4 #( .INIT(16'h7350) )  \n_response_1_1_iv_0_0[34]  (.A(
        \response[34]_net_1 ), .B(\response[33]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[34]_net_1 ));
    CFG4 #( .INIT(16'hBA98) )  \n_response_360_0[0]  (.A(m17_d_s), .B(
        m17_s), .C(m17_d_d), .D(i4_mux_0), .Y(
        \n_response_360_0[0]_net_1 ));
    SLE no_crc (.D(no_crc_397_net_1), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(no_crc_net_1));
    CFG3 #( .INIT(8'h80) )  \state_ns_0_a3_0_a2_0_a3[6]  (.A(
        \state_ns_0_a3_0_a2_0_a3_1[6]_net_1 ), .B(N_374), .C(N_393), 
        .Y(\state_ns[6] ));
    CFG3 #( .INIT(8'h80) )  un105_i_a3_0_0_RNIMG8H (.A(\arg[7]_net_1 ), 
        .B(N_3641), .C(\arg[6]_net_1 ), .Y(
        buffer_under_runlde_0_a6_0_1));
    CFG4 #( .INIT(16'h0010) )  un1_arg_12_3 (.A(\arg[4]_net_1 ), .B(
        \arg[5]_net_1 ), .C(\arg[27]_net_1 ), .D(\arg[6]_net_1 ), .Y(
        un1_arg_12_3_0));
    CFG4 #( .INIT(16'h7350) )  \n_response_1_1_iv_0_0[37]  (.A(
        \response[37]_net_1 ), .B(\response[36]_net_1 ), .C(N_3595), 
        .D(N_845), .Y(\n_response_1_1_iv_0_0[37]_net_1 ));
    CFG4 #( .INIT(16'h5551) )  \response_RNO[36]  (.A(
        \n_response_1_1_iv_0_0[36]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_response_1_sqmuxa_net_1), .D(n_state_0_sqmuxa), .Y(
        \n_response_1_1_iv_i[36] ));
    SLE crc_en (.D(N_3522_i), .CLK(sdclk_n_1), .EN(N_1699), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(crc_en_net_1));
    CFG3 #( .INIT(8'hFE) )  n_response_7_sqmuxa_1_0_0_o2 (.A(
        \arg[11]_net_1 ), .B(\arg[12]_net_1 ), .C(\arg[10]_net_1 ), .Y(
        N_229));
    CFG1 #( .INIT(2'h1) )  dsd_clkr_RNO (.A(dsd_clkr_net_1), .Y(
        dsd_clkr_i_i));
    CFG4 #( .INIT(16'h4000) )  un103_i_a6 (.A(N_3696), .B(N_3762), .C(
        N_1697), .D(un103_i_a6_0_net_1), .Y(un103_i_a6_net_1));
    CFG4 #( .INIT(16'h1000) )  \n_response_cnst_4_7_0_.m42_0_a3_1  (.A(
        \arg[14]_net_1 ), .B(\arg[13]_net_1 ), .C(\arg[9]_net_1 ), .D(
        N_372), .Y(N_335));
    CFG4 #( .INIT(16'h5070) )  response_ret_5_RNO (.A(
        \bus_state[3]_net_1 ), .B(N_202), .C(\n_response_406_m_0[11] ), 
        .D(N_3690), .Y(\n_response_406_m[11] ));
    CFG4 #( .INIT(16'hFFFE) )  \state_ns_0_i_o2[0]  (.A(
        \state_ns_0_i_o2_0[0]_net_1 ), .B(N_89), .C(
        \state_ns_0_i_o2_1[0]_net_1 ), .D(N_216), .Y(N_416));
    CFG2 #( .INIT(4'h2) )  n_cmd_out_iv_0_a2_9 (.A(\i[5]_net_1 ), .B(
        no_crc_net_1), .Y(N_174));
    CFG4 #( .INIT(16'hFFFE) )  \n_response_1_0_iv[0]  (.A(
        \n_response_49_m[0] ), .B(\n_response_1_0_iv_1[0]_net_1 ), .C(
        \n_response_360_m[0] ), .D(\n_response_123_m[0]_net_1 ), .Y(
        \n_response_1[0] ));
    CFG4 #( .INIT(16'h00CE) )  \state_RNO[9]  (.A(\state[6]_net_1 ), 
        .B(\state[9]_net_1 ), .C(N_221), .D(N_2221), .Y(N_2163_i));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNICPN85[4]  (.A(
        VCC_net_1), .B(\buffer_under_run[4]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[3] ), .S(\buffer_under_run_s[4] ), .Y(), 
        .FCO(\buffer_under_run_cry[4] ));
    SLE \response[31]  (.D(\n_response_1[31] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[31]_net_1 ));
    SLE response_ret_14 (.D(\response[8]_net_1 ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response_reto[8] ));
    CFG3 #( .INIT(8'hFB) )  \state_ns_0_o3[7]  (.A(\i[3] ), .B(N_276), 
        .C(\i[2] ), .Y(N_2181));
    CFG4 #( .INIT(16'h3A0A) )  i_cry_cy_424 (.A(\i_s_reto[0] ), .B(
        \i_reto[0] ), .C(N_3732_reto), .D(N_2431_reto), .Y(\i_0[0] ));
    CFG4 #( .INIT(16'hFFF8) )  \n_response_1_0_iv_2[3]  (.A(
        \state[12]_net_1 ), .B(\n_response_49[3]_net_1 ), .C(
        \n_response_159_m[3]_net_1 ), .D(
        \n_response_1_0_iv_0[3]_net_1 ), .Y(
        \n_response_1_0_iv_2[3]_net_1 ));
    CFG4 #( .INIT(16'hFEF0) )  \state_RNO[4]  (.A(un1_i_3), .B(
        n_crc_en_1_sqmuxa_i_o2_RNIVR871_net_1), .C(\state[3]_net_1 ), 
        .D(\state[4]_net_1 ), .Y(N_2223_i));
    CFG4 #( .INIT(16'hFFFE) )  \state_ns_0_i_o2_0[0]  (.A(N_216), .B(
        \state_ns_0_i_o2_0_3[0]_net_1 ), .C(N_360), .D(
        \state_ns_0_i_o2_0_0[0]_net_1 ), .Y(N_417));
    CFG4 #( .INIT(16'h0001) )  \state_ns_0_a3_0_a2_0_a3_1[6]  (.A(
        \bus_state[4]_net_1 ), .B(\ind[1]_net_1 ), .C(\ind[0]_net_1 ), 
        .D(\ind[3]_net_1 ), .Y(\state_ns_0_a3_0_a2_0_a3_1[6]_net_1 ));
    CFG4 #( .INIT(16'h3A0A) )  \i_lm_0[0]  (.A(\i_s_reto[0] ), .B(
        \i_reto[0] ), .C(N_3732_reto), .D(N_2431_reto), .Y(\i[0] ));
    CFG3 #( .INIT(8'h20) )  crc_en_RNO (.A(N_845), .B(N_3528), .C(
        N_244), .Y(N_3522_i));
    SLE \response[33]  (.D(\n_response_1[33] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[33]_net_1 ));
    SLE \i[4]  (.D(\i_lm[4] ), .CLK(sdclk_n_1), .EN(VCC_net_1), .ALn(
        u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    SLE \arg[2]  (.D(\n_arg[2]_net_1 ), .CLK(sdclk_n_1), .EN(un77), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\arg[2]_net_1 ));
    CFG4 #( .INIT(16'h7430) )  ind_394 (.A(\state[0]_net_1 ), .B(
        N_3524), .C(\ind[5]_net_1 ), .D(\ind[4]_net_1 ), .Y(
        ind_394_net_1));
    CFG4 #( .INIT(16'h0100) )  \arg_RNIDVHN1[4]  (.A(\arg[5]_net_1 ), 
        .B(\arg[4]_net_1 ), .C(\arg[6]_net_1 ), .D(
        un1_arg_13_i_i_a2_0_13_2), .Y(un1_arg_13_i_i_a2_0_13_4));
    CFG4 #( .INIT(16'hFCDC) )  \bus_state_ns_0[3]  (.A(
        \bus_state_ns_0_1[3]_net_1 ), .B(\bus_state_ns_0_0[3]_net_1 ), 
        .C(\bus_state[3]_net_1 ), .D(n_state_0_sqmuxa), .Y(
        \bus_state_ns[3] ));
    CFG4 #( .INIT(16'h3313) )  \state_RNO[1]  (.A(N_317_1), .B(
        \state_ns_i_0_0_0[1]_net_1 ), .C(\ind[3]_net_1 ), .D(
        \state[0]_net_1 ), .Y(N_2153_i));
    CFG4 #( .INIT(16'h0008) )  n_response_5_sqmuxa_1_1 (.A(
        \bus_state[3]_net_1 ), .B(N_1060), .C(\arg[26]_net_1 ), .D(
        \arg[27]_net_1 ), .Y(n_response_5_sqmuxa_1_1_net_1));
    CFG4 #( .INIT(16'h0010) )  \state_ns_0_a2_3_1_a6_0_a2_3[0]  (.A(
        \arg[26]_net_1 ), .B(\arg[17]_net_1 ), .C(\arg[16]_net_1 ), .D(
        N_221), .Y(\state_ns_0_a2_3_1_a6_0_a2_3[0]_net_1 ));
    SLE response_ret_8 (.D(\n_response_cnst_1_m[9] ), .CLK(sdclk_n_1), 
        .EN(un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \n_response_cnst_1_m_reto_0[9] ));
    CFG4 #( .INIT(16'hFFEC) )  \n_response_1_0_iv[2]  (.A(
        \state[9]_net_1 ), .B(\n_response_123_m[2]_net_1 ), .C(
        \n_response_360[2]_net_1 ), .D(\n_response_1_0_iv_2[2]_net_1 ), 
        .Y(\n_response_1[2] ));
    CFG4 #( .INIT(16'hFFF8) )  n_response_7_sqmuxa_1_0_0_tz_1 (.A(
        N_229), .B(\arg[13]_net_1 ), .C(N_10), .D(N_372), .Y(
        n_response_7_sqmuxa_1_0_0_tz_1_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \n_response_cnst_4_7_0_.m42_0_2  (.A(
        N_336), .B(N_335), .C(N_333), .D(N_337), .Y(m42_0_2));
    CFG2 #( .INIT(4'h8) )  \n_response_1_1_iv_0_a6_0[33]  (.A(N_845), 
        .B(\response[32]_net_1 ), .Y(N_3713));
    CFG2 #( .INIT(4'hD) )  n_response193_1_0_a3_0_o2 (.A(
        \arg[9]_net_1 ), .B(\arg[12]_net_1 ), .Y(N_3592));
    CFG3 #( .INIT(8'hAC) )  \n_response_cnst_4_7_0_.m6  (.A(N_702_1), 
        .B(N_4), .C(\arg[13]_net_1 ), .Y(i4_mux_0));
    CFG4 #( .INIT(16'h0008) )  n_response_16_sqmuxa_i_0_a3_1 (.A(
        \arg[13]_net_1 ), .B(\arg[11]_net_1 ), .C(N_4054), .D(N_4053), 
        .Y(N_313));
    CFG2 #( .INIT(4'h4) )  \n_arg_i_i_a3[0]  (.A(\state[0]_net_1 ), .B(
        cmd_q_net_1), .Y(N_342));
    CFG3 #( .INIT(8'h27) )  \n_response_1_0_iv_2_RNO_1[1]  (.A(N_706), 
        .B(\sound_card_ctrl[1]_net_1 ), .C(en49_c), .Y(
        \n_response_49_4_1_0[1] ));
    CFG4 #( .INIT(16'hAF3F) )  \n_i_iv_0[1]  (.A(\state[1]_net_1 ), .B(
        N_3589_i), .C(N_1696_i), .D(N_96_i), .Y(\n_i[1] ));
    CFG3 #( .INIT(8'h08) )  \bus_state_ns_0_a4_1_1[3]  (.A(
        \bus_state[2]_net_1 ), .B(\state[0]_net_1 ), .C(data_bus_busy), 
        .Y(\bus_state_ns_0_a4_1_1[3]_net_1 ));
    CFG4 #( .INIT(16'h0ACC) )  arg_366 (.A(\arg[20]_net_1 ), .B(
        \arg[21]_net_1 ), .C(\state[0]_net_1 ), .D(un77), .Y(
        arg_366_net_1));
    CFG2 #( .INIT(4'h8) )  un12_n_i_ac0_5 (.A(un12_n_i_c3), .B(\i[3] ), 
        .Y(un12_n_i_c4));
    SLE \state[9]  (.D(N_2163_i), .CLK(sdclk_n_1), .EN(VCC_net_1), 
        .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[9]_net_1 ));
    CFG4 #( .INIT(16'hFF0E) )  un96_i_0 (.A(\state[4]_net_1 ), .B(
        \state[0]_net_1 ), .C(\state[1]_net_1 ), .D(N_3745), .Y(
        un96_i_0_net_1));
    CFG3 #( .INIT(8'hEA) )  \n_response_1_1_iv_0[24]  (.A(
        \n_response_1_1_iv_0_0[24]_net_1 ), .B(un1_n_bit_0_sqmuxa_i_0), 
        .C(n_state_1_sqmuxa), .Y(\n_response_1[24] ));
    CFG2 #( .INIT(4'h9) )  \i_qxu[0]  (.A(N_845), .B(\i[0] ), .Y(
        \i_qxu[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \n_response_36_0[7]  (.A(N_1163), .B(
        \buffer_under_run[7]_net_1 ), .Y(N_2541));
    CFG4 #( .INIT(16'h88A0) )  \n_response_1_0_iv_RNO_0[0]  (.A(
        \state[9]_net_1 ), .B(\response[0]_net_1 ), .C(
        \n_response_360_1[0]_net_1 ), .D(N_709), .Y(
        \n_response_360_m[0] ));
    SLE \response[14]  (.D(\n_response_1[14] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[14]_net_1 ));
    SLE \response[24]  (.D(\n_response_1[24] ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \response[24]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \buffer_under_run_RNIG4NC2[1]  (.A(
        VCC_net_1), .B(\buffer_under_run[1]_net_1 ), .C(
        \state[12]_net_1 ), .D(GND_net_1), .FCI(
        \buffer_under_run_cry[0] ), .S(\buffer_under_run_s[1] ), .Y(), 
        .FCO(\buffer_under_run_cry[1] ));
    CFG4 #( .INIT(16'h4447) )  \n_response_1_0_iv_2_RNO_2[1]  (.A(
        \response[1] ), .B(\arg[31]_net_1 ), .C(N_702), .D(N_706), .Y(
        \n_response_49_4_1_1[1] ));
    CFG3 #( .INIT(8'hFE) )  \bus_state_ns_0_o3_0[3]  (.A(
        \state[10]_net_1 ), .B(n_state_0_sqmuxa), .C(N_1686_i), .Y(
        N_2265));
    SLE response_ret_3 (.D(\state[9]_net_1 ), .CLK(sdclk_n_1), .EN(
        un1_state_11_i), .ALn(u8_sb_0_HPMS_READY), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_reto[9] ));
    CFG3 #( .INIT(8'hA8) )  \bus_state_ns_0_0_a2[1]  (.A(
        \bus_state[1]_net_1 ), .B(N_2266), .C(N_2265), .Y(N_3624));
    CFG4 #( .INIT(16'h3732) )  \n_response_49[6]  (.A(\arg[31]_net_1 ), 
        .B(\n_response_49_1_1[6]_net_1 ), .C(N_702), .D(
        \n_response_36[6]_net_1 ), .Y(\n_response_49[6]_net_1 ));
    CFG4 #( .INIT(16'hF700) )  un1_buffer_under_runlto5_RNI8UTG2 (.A(
        \buffer_under_run[7]_net_1 ), .B(\buffer_under_run[6]_net_1 ), 
        .C(un1_buffer_under_runlt7), .D(buffer_under_runlde_0_a6_5), 
        .Y(buffer_under_runlde_0_a6_7));
    CFG4 #( .INIT(16'h2000) )  \state_ns_0_a3_0_a2_0_a3_4[2]  (.A(
        \i[5]_net_1 ), .B(\i[4]_net_1 ), .C(\i[0] ), .D(\i[3] ), .Y(
        N_318_4));
    CFG4 #( .INIT(16'hAE0C) )  \n_response_1_0_iv_0[9]  (.A(
        \response[9] ), .B(\state[10]_net_1 ), .C(N_1060), .D(N_3595), 
        .Y(\n_response_1_0_iv_0[9]_net_1 ));
    
endmodule


module clock138master(
       reset_n_i,
       en45_c,
       en49_c,
       u8_sb_0_HPMS_READY,
       clock138_data_c,
       clock138_lrck_c,
       clock138_bck_c,
       reset_n_i_i
    );
output reset_n_i;
input  en45_c;
input  en49_c;
input  u8_sb_0_HPMS_READY;
output clock138_data_c;
input  clock138_lrck_c;
input  clock138_bck_c;
input  reset_n_i_i;

    wire \i[0]_net_1 , \i_s[0] , work_net_1, VCC_net_1, n_work4_net_1, 
        GND_net_1, olrck_net_1, i4_mux, n_i6_net_1, \i[1]_net_1 , 
        \i_s[1] , \i[2]_net_1 , \i_s[2] , \i[3]_net_1 , \i_s[3] , 
        \i[4]_net_1 , \i_s[4] , \i[5]_net_1 , \i_s[5] , \i[6]_net_1 , 
        \i_s[6] , \i[7]_net_1 , \i_s[7] , \i[8]_net_1 , \i_s[8] , 
        \i[9]_net_1 , \i_s[9] , \i[10]_net_1 , \i_s[10] , 
        \i[11]_net_1 , \i_s[11] , \i[12]_net_1 , \i_s[12] , 
        \i[13]_net_1 , \i_s[13] , \i[14]_net_1 , \i_s[14]_net_1 , 
        i_s_412_FCO, \i_cry[1]_net_1 , \i_cry[2]_net_1 , 
        \i_cry[3]_net_1 , \i_cry[4]_net_1 , \i_cry[5]_net_1 , 
        \i_cry[6]_net_1 , \i_cry[7]_net_1 , \i_cry[8]_net_1 , 
        \i_cry[9]_net_1 , \i_cry[10]_net_1 , \i_cry[11]_net_1 , 
        \i_cry[12]_net_1 , \i_cry[13]_net_1 , m10_am_1, m5, m10_am, 
        m10_bm, m7;
    
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[12]  (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[11]_net_1 ), .S(\i_s[12] ), .Y(), .FCO(
        \i_cry[12]_net_1 ));
    CFG3 #( .INIT(8'hA8) )  reset_n_i_inst_1 (.A(u8_sb_0_HPMS_READY), 
        .B(en49_c), .C(en45_c), .Y(reset_n_i));
    SLE work (.D(VCC_net_1), .CLK(clock138_bck_c), .EN(n_work4_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(work_net_1));
    SLE \i[9]  (.D(\i_s[9] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    SLE \i[2]  (.D(\i_s[2] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[10]  (.D(\i_s[10] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[10]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  i_s_412 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(i_s_412_FCO));
    SLE \i[3]  (.D(\i_s[3] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    SLE \i[8]  (.D(\i_s[8] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h8D) )  \key_pmux_0_0_0_.m10_am  (.A(\i[9]_net_1 ), 
        .B(m5), .C(m10_am_1), .Y(m10_am));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[8]  (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[7]_net_1 ), .S(\i_s[8] ), .Y(), .FCO(\i_cry[8]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \key_pmux_0_0_0_.m10_ns  (.A(m10_bm), .B(
        \i[12]_net_1 ), .C(m10_am), .Y(i4_mux));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(\i_cry[5]_net_1 ));
    CFG2 #( .INIT(4'h9) )  \key_pmux_0_0_0_.m5  (.A(\i[7]_net_1 ), .B(
        \i[10]_net_1 ), .Y(m5));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(i_s_412_FCO), 
        .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG1 #( .INIT(2'h1) )  \i_RNO[0]  (.A(\i[0]_net_1 ), .Y(\i_s[0] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[11]  (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[10]_net_1 ), .S(\i_s[11] ), .Y(), .FCO(
        \i_cry[11]_net_1 ));
    SLE \i[14]  (.D(\i_s[14]_net_1 ), .CLK(clock138_bck_c), .EN(
        n_i6_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[14]_net_1 ));
    SLE \i[0]  (.D(\i_s[0] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    CFG2 #( .INIT(4'h2) )  n_work4 (.A(olrck_net_1), .B(
        clock138_lrck_c), .Y(n_work4_net_1));
    SLE \i[13]  (.D(\i_s[13] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[13]_net_1 ));
    CFG4 #( .INIT(16'hB3C4) )  \key_pmux_0_0_0_.m10_bm  (.A(
        \i[11]_net_1 ), .B(\i[9]_net_1 ), .C(m7), .D(m5), .Y(m10_bm));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[9]  (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[8]_net_1 ), .S(\i_s[9] ), .Y(), .FCO(\i_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[13]  (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[12]_net_1 ), .S(\i_s[13] ), .Y(), .FCO(
        \i_cry[13]_net_1 ));
    SLE \i[5]  (.D(\i_s[5] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \key_pmux_0_0_0_.m7  (.A(\i[7]_net_1 ), .B(
        \i[10]_net_1 ), .Y(m7));
    SLE olrck (.D(clock138_lrck_c), .CLK(clock138_bck_c), .EN(
        VCC_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(olrck_net_1));
    SLE \i[6]  (.D(\i_s[6] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    SLE \i[12]  (.D(\i_s[12] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[10]  (.A(VCC_net_1), .B(
        \i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[9]_net_1 ), .S(\i_s[10] ), .Y(), .FCO(\i_cry[10]_net_1 )
        );
    CFG3 #( .INIT(8'h2A) )  n_i6 (.A(work_net_1), .B(\i[14]_net_1 ), 
        .C(\i[13]_net_1 ), .Y(n_i6_net_1));
    SLE key_pmux_0_dreg (.D(i4_mux), .CLK(clock138_bck_c), .EN(
        n_i6_net_1), .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clock138_data_c));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    SLE \i[7]  (.D(\i_s[7] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    SLE \i[4]  (.D(\i_s[4] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    CFG4 #( .INIT(16'h2ABB) )  \key_pmux_0_0_0_.m10_am_1  (.A(
        \i[7]_net_1 ), .B(\i[10]_net_1 ), .C(\i[8]_net_1 ), .D(
        \i[11]_net_1 ), .Y(m10_am_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_s[14]  (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[13]_net_1 ), .S(\i_s[14]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(\i_cry[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[6]_net_1 ), .S(\i_s[7] ), .Y(), .FCO(\i_cry[7]_net_1 ));
    SLE \i[1]  (.D(\i_s[1] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    SLE \i[11]  (.D(\i_s[11] ), .CLK(clock138_bck_c), .EN(n_i6_net_1), 
        .ALn(reset_n_i_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[11]_net_1 ));
    
endmodule


module test(
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0,
       test_0_HWDATA,
       test_0_HADDR,
       test_0_HADDR_i_0,
       test_0_HTRANS_0,
       reset_n_i_i_3,
       clock138_bck_c,
       clock138_lrck_c,
       clock138_data_c,
       reset_n_i,
       u8_sb_0_HPMS_READY,
       en45_c,
       en49_c,
       spdif_en_c,
       reset_n_i_i_2,
       reset_n_i_0,
       reset_n_i_i_1,
       reset_n_i_1,
       reset_n_i_i_0,
       reset_n_i_3,
       reset_n_i_i,
       reset_n_i_2,
       spdif_tx_c,
       test_0_HWRITE,
       u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0,
       mclk_c,
       cmd,
       sd_d0,
       sd_d1,
       sd_d2,
       sd_d3,
       obck,
       olrck,
       odata,
       sdclk_c
    );
input  [31:0] u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0;
output [31:0] test_0_HWDATA;
output [16:2] test_0_HADDR;
output test_0_HADDR_i_0;
output test_0_HTRANS_0;
input  reset_n_i_i_3;
input  clock138_bck_c;
input  clock138_lrck_c;
output clock138_data_c;
output reset_n_i;
input  u8_sb_0_HPMS_READY;
output en45_c;
output en49_c;
output spdif_en_c;
input  reset_n_i_i_2;
output reset_n_i_0;
input  reset_n_i_i_1;
output reset_n_i_1;
input  reset_n_i_i_0;
output reset_n_i_3;
input  reset_n_i_i;
output reset_n_i_2;
output spdif_tx_c;
output test_0_HWRITE;
input  u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0;
input  mclk_c;
inout  cmd;
inout  sd_d0;
inout  sd_d1;
inout  sd_d2;
inout  sd_d3;
inout  obck;
inout  olrck;
inout  odata;
input  sdclk_c;

    wire sdclk_n_1, sdclk_n_i, sdclk_c_i, odata_i, odata_o, VCC_net_1, 
        olrck_i, olrck_o, obck_i, obck_o, \sd_data_in[3] , 
        \sd_data_out[3] , sd_data_out_en_i_i, \sd_data_in[2] , 
        \sd_data_out[2] , \sd_data_in[1] , \sd_data_out[1] , 
        data_out_en_ret_fast_i, \sd_data_in[0] , \sd_data_out[0] , 
        cmd_in, cmd_out, cmd_out_en_i_i, mclk_1, GND_net_1;
    
    BIBUF UDAT22 (.PAD(odata), .D(odata_o), .E(VCC_net_1), .Y(odata_i));
    CFG1 #( .INIT(2'h1) )  UCK3_RNO (.A(sdclk_c), .Y(sdclk_c_i));
    GND GND (.Y(GND_net_1));
    CLKINT_PRESERVE UCK3 (.A(sdclk_c_i), .Y(sdclk_n_1));
    BIBUF UDAT2 (.PAD(sd_d2), .D(\sd_data_out[2] ), .E(
        sd_data_out_en_i_i), .Y(\sd_data_in[2] ));
    BIBUF UDAT1 (.PAD(sd_d1), .D(\sd_data_out[1] ), .E(
        data_out_en_ret_fast_i), .Y(\sd_data_in[1] ));
    BIBUF UBB (.PAD(cmd), .D(cmd_out), .E(cmd_out_en_i_i), .Y(cmd_in));
    sdtop u100 (.test_0_HADDR({test_0_HADDR[16], test_0_HADDR[15], 
        test_0_HADDR[14], test_0_HADDR[13], test_0_HADDR[12], 
        test_0_HADDR[11], test_0_HADDR[10], test_0_HADDR[9], 
        test_0_HADDR[8], test_0_HADDR[7], test_0_HADDR[6], 
        test_0_HADDR[5], test_0_HADDR[4], test_0_HADDR[3], 
        test_0_HADDR[2]}), .test_0_HWDATA({test_0_HWDATA[31], 
        test_0_HWDATA[30], test_0_HWDATA[29], test_0_HWDATA[28], 
        test_0_HWDATA[27], test_0_HWDATA[26], test_0_HWDATA[25], 
        test_0_HWDATA[24], test_0_HWDATA[23], test_0_HWDATA[22], 
        test_0_HWDATA[21], test_0_HWDATA[20], test_0_HWDATA[19], 
        test_0_HWDATA[18], test_0_HWDATA[17], test_0_HWDATA[16], 
        test_0_HWDATA[15], test_0_HWDATA[14], test_0_HWDATA[13], 
        test_0_HWDATA[12], test_0_HWDATA[11], test_0_HWDATA[10], 
        test_0_HWDATA[9], test_0_HWDATA[8], test_0_HWDATA[7], 
        test_0_HWDATA[6], test_0_HWDATA[5], test_0_HWDATA[4], 
        test_0_HWDATA[3], test_0_HWDATA[2], test_0_HWDATA[1], 
        test_0_HWDATA[0]}), .u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0({
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1], 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0]}), .sd_data_in({
        \sd_data_in[3] , \sd_data_in[2] , \sd_data_in[1] , 
        \sd_data_in[0] }), .sd_data_out({\sd_data_out[3] , 
        \sd_data_out[2] , \sd_data_out[1] , \sd_data_out[0] }), 
        .test_0_HTRANS_0(test_0_HTRANS_0), .test_0_HADDR_i_0(
        test_0_HADDR_i_0), .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .test_0_HWRITE(
        test_0_HWRITE), .spdif_tx_c(spdif_tx_c), .olrck_o(olrck_o), 
        .reset_n_i_2(reset_n_i_2), .reset_n_i_i_2(reset_n_i_i), 
        .reset_n_i_3(reset_n_i_3), .reset_n_i_i_1(reset_n_i_i_0), 
        .reset_n_i_1(reset_n_i_1), .reset_n_i_i_0(reset_n_i_i_1), 
        .reset_n_i_0(reset_n_i_0), .mclk_1(mclk_1), .reset_n_i_i(
        reset_n_i_i_2), .sd_data_out_en_i_i(sd_data_out_en_i_i), 
        .data_out_en_ret_fast_i(data_out_en_ret_fast_i), .odata_o(
        odata_o), .obck_o(obck_o), .cmd_in(cmd_in), .sdclk_n_i(
        sdclk_n_i), .cmd_out(cmd_out), .spdif_en_c(spdif_en_c), 
        .en49_c(en49_c), .en45_c(en45_c), .sdclk_n_1(sdclk_n_1), 
        .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY), .cmd_out_en_i_i(
        cmd_out_en_i_i));
    VCC VCC (.Y(VCC_net_1));
    BIBUF UDAT3 (.PAD(sd_d3), .D(\sd_data_out[3] ), .E(
        sd_data_out_en_i_i), .Y(\sd_data_in[3] ));
    CLKINT_PRESERVE UCK1 (.A(mclk_c), .Y(mclk_1));
    BIBUF UDAT0 (.PAD(sd_d0), .D(\sd_data_out[0] ), .E(
        data_out_en_ret_fast_i), .Y(\sd_data_in[0] ));
    BIBUF UDAT21 (.PAD(olrck), .D(olrck_o), .E(VCC_net_1), .Y(olrck_i));
    clock138master u200 (.reset_n_i(reset_n_i), .en45_c(en45_c), 
        .en49_c(en49_c), .u8_sb_0_HPMS_READY(u8_sb_0_HPMS_READY), 
        .clock138_data_c(clock138_data_c), .clock138_lrck_c(
        clock138_lrck_c), .clock138_bck_c(clock138_bck_c), 
        .reset_n_i_i(reset_n_i_i_3));
    CFG1 #( .INIT(2'h1) )  UCK3_RNIJ7S9 (.A(sdclk_n_1), .Y(sdclk_n_i));
    BIBUF UDAT20 (.PAD(obck), .D(obck_o), .E(VCC_net_1), .Y(obck_i));
    
endmodule


module u8(
       DEVRST_N,
       clock138_bck,
       clock138_lrck,
       mclk,
       sdclk,
       clock138_data,
       en45,
       en49,
       led0,
       led1,
       led2,
       led3,
       led4,
       led5,
       led6,
       led7,
       sd_det,
       spdif_en,
       spdif_tx,
       cmd,
       obck,
       odata,
       olrck,
       sd_d0,
       sd_d1,
       sd_d2,
       sd_d3
    );
input  DEVRST_N;
input  clock138_bck;
input  clock138_lrck;
input  mclk;
input  sdclk;
output clock138_data;
output en45;
output en49;
output led0;
output led1;
output led2;
output led3;
output led4;
output led5;
output led6;
output led7;
output sd_det;
output spdif_en;
output spdif_tx;
inout  cmd;
inout  obck;
inout  odata;
inout  olrck;
inout  sd_d0;
inout  sd_d1;
inout  sd_d2;
inout  sd_d3;

    wire u8_sb_0_HPMS_READY, \test_0_HADDR[15] , \test_0_HADDR[16] , 
        \test_0_HTRANS[1] , test_0_HWRITE, \test_0_HWDATA[0] , 
        \test_0_HWDATA[1] , \test_0_HWDATA[2] , \test_0_HWDATA[3] , 
        \test_0_HWDATA[4] , \test_0_HWDATA[5] , \test_0_HWDATA[6] , 
        \test_0_HWDATA[7] , \test_0_HWDATA[8] , \test_0_HWDATA[9] , 
        \test_0_HWDATA[10] , \test_0_HWDATA[11] , \test_0_HWDATA[12] , 
        \test_0_HWDATA[13] , \test_0_HWDATA[14] , \test_0_HWDATA[15] , 
        \test_0_HWDATA[16] , \test_0_HWDATA[17] , \test_0_HWDATA[18] , 
        \test_0_HWDATA[19] , \test_0_HWDATA[20] , \test_0_HWDATA[21] , 
        \test_0_HWDATA[22] , \test_0_HWDATA[23] , \test_0_HWDATA[24] , 
        \test_0_HWDATA[25] , \test_0_HWDATA[26] , \test_0_HWDATA[27] , 
        \test_0_HWDATA[28] , \test_0_HWDATA[29] , \test_0_HWDATA[30] , 
        \test_0_HWDATA[31] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31] , 
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0, VCC_net_1, GND_net_1, 
        clock138_bck_c, clock138_lrck_c, mclk_c, sdclk_c, 
        clock138_data_c, en45_c, en49_c, spdif_en_c, spdif_tx_c, 
        \test_0_HADDR[14] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10] , 
        \test_0_HADDR[2] , \test_0_HADDR[3] , \test_0_HADDR[4] , 
        \test_0_HADDR[5] , \test_0_HADDR[6] , \test_0_HADDR[7] , 
        \test_0_HADDR[8] , \test_0_HADDR[9] , \test_0_HADDR[10] , 
        \test_0_HADDR[11] , \test_0_HADDR[12] , \test_0_HADDR[13] , 
        \test_0_HADDR_i[16] , \test_0.u200.reset_n_i_i , 
        \test_0.u100.USPDIF_TX.reset_n_i_i , 
        \test_0.u100.UPCMTX.reset_n_i_i , 
        \test_0.u100.UDOP.reset_n_i_i , 
        \test_0.u100.UDSDTX.reset_n_i_i , reset_n_i_3, reset_n_i_2, 
        reset_n_i_1, reset_n_i_0, reset_n_i, clock138_bck_ibuf_net_1;
    
    OUTBUF clock138_data_obuf (.D(clock138_data_c), .PAD(clock138_data)
        );
    OUTBUF spdif_en_obuf (.D(spdif_en_c), .PAD(spdif_en));
    TRIBUFF led4_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(led4));
    u8_sb u8_sb_0 (.u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0({
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0] }), 
        .test_0_HWDATA({\test_0_HWDATA[31] , \test_0_HWDATA[30] , 
        \test_0_HWDATA[29] , \test_0_HWDATA[28] , \test_0_HWDATA[27] , 
        \test_0_HWDATA[26] , \test_0_HWDATA[25] , \test_0_HWDATA[24] , 
        \test_0_HWDATA[23] , \test_0_HWDATA[22] , \test_0_HWDATA[21] , 
        \test_0_HWDATA[20] , \test_0_HWDATA[19] , \test_0_HWDATA[18] , 
        \test_0_HWDATA[17] , \test_0_HWDATA[16] , \test_0_HWDATA[15] , 
        \test_0_HWDATA[14] , \test_0_HWDATA[13] , \test_0_HWDATA[12] , 
        \test_0_HWDATA[11] , \test_0_HWDATA[10] , \test_0_HWDATA[9] , 
        \test_0_HWDATA[8] , \test_0_HWDATA[7] , \test_0_HWDATA[6] , 
        \test_0_HWDATA[5] , \test_0_HWDATA[4] , \test_0_HWDATA[3] , 
        \test_0_HWDATA[2] , \test_0_HWDATA[1] , \test_0_HWDATA[0] }), 
        .test_0_HADDR({\test_0_HADDR[16] , \test_0_HADDR[15] , 
        \test_0_HADDR[14] , \test_0_HADDR[13] , \test_0_HADDR[12] , 
        \test_0_HADDR[11] , \test_0_HADDR[10] , \test_0_HADDR[9] , 
        \test_0_HADDR[8] , \test_0_HADDR[7] , \test_0_HADDR[6] , 
        \test_0_HADDR[5] , \test_0_HADDR[4] , \test_0_HADDR[3] , 
        \test_0_HADDR[2] }), .test_0_HADDR_i_0(\test_0_HADDR_i[16] ), 
        .test_0_HTRANS_0(\test_0_HTRANS[1] ), .u8_sb_0_HPMS_READY(
        u8_sb_0_HPMS_READY), .test_0_HWRITE(test_0_HWRITE), 
        .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .mclk_c(mclk_c), 
        .DEVRST_N(DEVRST_N));
    CLKINT clock138_bck_ibuf_RNIS2E8 (.A(clock138_bck_ibuf_net_1), .Y(
        clock138_bck_c));
    INBUF mclk_ibuf (.PAD(mclk), .Y(mclk_c));
    OUTBUF spdif_tx_obuf (.D(spdif_tx_c), .PAD(spdif_tx));
    GND GND (.Y(GND_net_1));
    OUTBUF led1_obuf (.D(GND_net_1), .PAD(led1));
    CLKINT I_431 (.A(reset_n_i_0), .Y(\test_0.u100.UDSDTX.reset_n_i_i )
        );
    CLKINT I_434 (.A(reset_n_i), .Y(\test_0.u200.reset_n_i_i ));
    OUTBUF en45_obuf (.D(en45_c), .PAD(en45));
    INBUF clock138_lrck_ibuf (.PAD(clock138_lrck), .Y(clock138_lrck_c));
    CLKINT I_430 (.A(reset_n_i_1), .Y(\test_0.u100.UPCMTX.reset_n_i_i )
        );
    test test_0 (.u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0({
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[31] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[30] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[29] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[28] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[27] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[26] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[25] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[24] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[23] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[22] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[21] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[20] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[19] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[18] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[17] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[16] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[15] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[14] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[13] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[12] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[11] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[10] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[9] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[8] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[7] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[6] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[5] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[4] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[3] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[2] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[1] , 
        \u8_sb_0_HPMS_FIC_0_USER_MASTER_HRDATA_M0[0] }), 
        .test_0_HWDATA({\test_0_HWDATA[31] , \test_0_HWDATA[30] , 
        \test_0_HWDATA[29] , \test_0_HWDATA[28] , \test_0_HWDATA[27] , 
        \test_0_HWDATA[26] , \test_0_HWDATA[25] , \test_0_HWDATA[24] , 
        \test_0_HWDATA[23] , \test_0_HWDATA[22] , \test_0_HWDATA[21] , 
        \test_0_HWDATA[20] , \test_0_HWDATA[19] , \test_0_HWDATA[18] , 
        \test_0_HWDATA[17] , \test_0_HWDATA[16] , \test_0_HWDATA[15] , 
        \test_0_HWDATA[14] , \test_0_HWDATA[13] , \test_0_HWDATA[12] , 
        \test_0_HWDATA[11] , \test_0_HWDATA[10] , \test_0_HWDATA[9] , 
        \test_0_HWDATA[8] , \test_0_HWDATA[7] , \test_0_HWDATA[6] , 
        \test_0_HWDATA[5] , \test_0_HWDATA[4] , \test_0_HWDATA[3] , 
        \test_0_HWDATA[2] , \test_0_HWDATA[1] , \test_0_HWDATA[0] }), 
        .test_0_HADDR({\test_0_HADDR[16] , \test_0_HADDR[15] , 
        \test_0_HADDR[14] , \test_0_HADDR[13] , \test_0_HADDR[12] , 
        \test_0_HADDR[11] , \test_0_HADDR[10] , \test_0_HADDR[9] , 
        \test_0_HADDR[8] , \test_0_HADDR[7] , \test_0_HADDR[6] , 
        \test_0_HADDR[5] , \test_0_HADDR[4] , \test_0_HADDR[3] , 
        \test_0_HADDR[2] }), .test_0_HADDR_i_0(\test_0_HADDR_i[16] ), 
        .test_0_HTRANS_0(\test_0_HTRANS[1] ), .reset_n_i_i_3(
        \test_0.u200.reset_n_i_i ), .clock138_bck_c(clock138_bck_c), 
        .clock138_lrck_c(clock138_lrck_c), .clock138_data_c(
        clock138_data_c), .reset_n_i(reset_n_i), .u8_sb_0_HPMS_READY(
        u8_sb_0_HPMS_READY), .en45_c(en45_c), .en49_c(en49_c), 
        .spdif_en_c(spdif_en_c), .reset_n_i_i_2(
        \test_0.u100.USPDIF_TX.reset_n_i_i ), .reset_n_i_0(reset_n_i_0)
        , .reset_n_i_i_1(\test_0.u100.UDSDTX.reset_n_i_i ), 
        .reset_n_i_1(reset_n_i_1), .reset_n_i_i_0(
        \test_0.u100.UPCMTX.reset_n_i_i ), .reset_n_i_3(reset_n_i_3), 
        .reset_n_i_i(\test_0.u100.UDOP.reset_n_i_i ), .reset_n_i_2(
        reset_n_i_2), .spdif_tx_c(spdif_tx_c), .test_0_HWRITE(
        test_0_HWRITE), .u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0(
        u8_sb_0_HPMS_FIC_0_USER_MASTER_HREADY_M0), .mclk_c(mclk_c), 
        .cmd(cmd), .sd_d0(sd_d0), .sd_d1(sd_d1), .sd_d2(sd_d2), .sd_d3(
        sd_d3), .obck(obck), .olrck(olrck), .odata(odata), .sdclk_c(
        sdclk_c));
    OUTBUF led2_obuf (.D(GND_net_1), .PAD(led2));
    CLKINT I_427 (.A(reset_n_i_3), .Y(\test_0.u100.UDOP.reset_n_i_i ));
    OUTBUF en49_obuf (.D(en49_c), .PAD(en49));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF sd_det_obuf (.D(GND_net_1), .PAD(sd_det));
    INBUF clock138_bck_ibuf (.PAD(clock138_bck), .Y(
        clock138_bck_ibuf_net_1));
    TRIBUFF led7_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(led7));
    OUTBUF led0_obuf (.D(GND_net_1), .PAD(led0));
    OUTBUF led3_obuf (.D(GND_net_1), .PAD(led3));
    CLKINT I_429 (.A(reset_n_i_2), .Y(
        \test_0.u100.USPDIF_TX.reset_n_i_i ));
    INBUF sdclk_ibuf (.PAD(sdclk), .Y(sdclk_c));
    TRIBUFF led6_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(led6));
    TRIBUFF led5_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(led5));
    
endmodule
